// Copyright 2022 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.
//

/*
 TODO_1: substitute the current ram_2p.sv for data and instr with the actuale sram_ctrl
 ip present in the opentitan repo (and change also the memory mapping for it, accordingly
 to the memory map used in opentitan).
 TODO_3: since the simulator control is not an opentitan ip, it could be possible to
 remove it and use the uart to print out the output of test softwares
*/

`include "prim_assert.sv"
`include "../../ip/tlul2axi/test/tlul_assign.svh"
`include "../../../../../deps/axi_scmi_mailbox/include/axi_typedef.svh"
`include "../../../../../deps/axi_scmi_mailbox/include/axi_assign.svh"

`ifndef RV32M
  `define RV32M ibex_pkg::RV32MFast
`endif

`ifndef RV32B
  `define RV32B ibex_pkg::RV32BNone
`endif

`ifndef RegFile
  `define RegFile ibex_pkg::RegFileFF
`endif


module opentitan 
  import axi_pkg::*;
  import jtag_pkg::*;
  #(

  // Manually defined parameters

  // Auto-inferred parameters
  // parameters for uart0
  // parameters for uart1
  // parameters for uart2
  // parameters for uart3
  // parameters for gpio
  // parameters for spi_device
  // parameters for spi_host0
  // parameters for spi_host1
  // parameters for i2c0
  // parameters for i2c1
  // parameters for i2c2
  // parameters for pattgen
  // parameters for rv_timer
  // parameters for usbdev
  // parameters for otp_ctrl
  parameter OtpCtrlMemInitFile = "/home/mciani/Workspace/cva6/hardware/working_dir/opentitan/hw/top_titangrey/examples/sw/simple_system/hello_test/otp-img.vmem",
  // parameters for lc_ctrl
  // parameters for alert_handler
  // parameters for pwrmgr_aon
  // parameters for rstmgr_aon
  // parameters for clkmgr_aon
  // parameters for sysrst_ctrl_aon
  // parameters for adc_ctrl_aon
  // parameters for pwm_aon
  // parameters for pinmux_aon
  parameter pinmux_pkg::target_cfg_t PinmuxAonTargetCfg = pinmux_pkg::DefaultTargetCfg,
  // parameters for aon_timer_aon
  // parameters for sensor_ctrl_aon
  // parameters for sram_ctrl_ret_aon
  parameter bit SramCtrlRetAonInstrExec = 0,
  // parameters for flash_ctrl
  // parameters for rv_dm
  parameter logic [31:0] RvDmIdcodeValue = 32'h 0000_0001,
  // parameters for rv_plic
  // parameters for aes
  parameter bit AesMasking = 1,
  parameter aes_pkg::sbox_impl_e AesSBoxImpl = aes_pkg::SBoxImplDom,
  parameter int unsigned SecAesStartTriggerDelay = 0,
  parameter bit SecAesAllowForcingMasks = 1'b0,
  parameter bit SecAesSkipPRNGReseeding = 1'b0,
  // parameters for hmac
  // parameters for kmac
  parameter bit KmacEnMasking = 1'b0, //1,
  parameter int KmacReuseShare = 0,
  // parameters for keymgr
  parameter bit KeymgrKmacEnMasking = 1'b0,//1,
  // parameters for csrng
  parameter aes_pkg::sbox_impl_e CsrngSBoxImpl = aes_pkg::SBoxImplCanright,
  // parameters for entropy_src
  parameter bit EntropySrcStub = 0,
  // parameters for edn0
  // parameters for edn1
  // parameters for sram_ctrl_main
  parameter bit SramCtrlMainInstrExec = 1,
  // parameters for otbn
  parameter bit OtbnStub = 0,
  parameter otbn_pkg::regfile_e OtbnRegFile = otbn_pkg::RegFileFF,
  // parameters for rom_ctrl
  parameter SRAMInitFile = "",//home/mciani/Workspace/cva6/hardware/working_dir/opentitan/hw/top_titangrey/examples/sw/simple_system/hello_test/ram.vmem",
  parameter RomCtrlBootRomInitFile = "/home/mciani/Workspace/cva6/hardware/working_dir/opentitan/hw/top_titangrey/examples/sw/simple_system/hello_test/scr_bootrom.vmem",
  parameter bit SecRomCtrlDisableScrambling = 1'b0,//1'b0,  
  // parameters for rv_core_ibex
  parameter bit RvCoreIbexPMPEnable = 0,//1
  parameter int unsigned RvCoreIbexPMPGranularity = 0,
  parameter int unsigned RvCoreIbexPMPNumRegions = 16,
  parameter int unsigned RvCoreIbexMHPMCounterNum = 10,
  parameter int unsigned RvCoreIbexMHPMCounterWidth = 32,
  parameter bit RvCoreIbexRV32E = 0,
  parameter ibex_pkg::rv32m_e RvCoreIbexRV32M = ibex_pkg::RV32MSingleCycle,
  parameter ibex_pkg::rv32b_e RvCoreIbexRV32B = ibex_pkg::RV32BNone,
  parameter ibex_pkg::regfile_e RvCoreIbexRegFile = ibex_pkg::RegFileFF,
  parameter bit RvCoreIbexBranchTargetALU = 1,
  parameter bit RvCoreIbexWritebackStage =1,
  parameter bit RvCoreIbexICache = 1,
  parameter bit RvCoreIbexICacheECC = 1,
  parameter bit RvCoreIbexBranchPredictor = 0,
  parameter bit RvCoreIbexDbgTriggerEn = 1,
  parameter bit RvCoreIbexSecureIbex = 1,
  parameter int unsigned RvCoreIbexDmHaltAddr =
      tl_main_pkg::ADDR_SPACE_RV_DM__ROM + dm::HaltAddress[31:0],
  parameter int unsigned RvCoreIbexDmExceptionAddr =
      tl_main_pkg::ADDR_SPACE_RV_DM__ROM + dm::ExceptionAddress[31:0],
  parameter bit RvCoreIbexPipeLine = 0,
  parameter type axi_req_t  = logic,
  parameter type axi_resp_t = logic
) (
  
  // spi_device
  input logic        cio_spi_device_sck_p2d,
  input logic        cio_spi_device_csb_p2d,
  input logic [3:0]  cio_spi_device_sd_p2d,
  output logic [3:0] cio_spi_device_sd_d2p,
  output logic [3:0] cio_spi_device_sd_en_d2p,
  // spi_host0
  input logic [3:0]  cio_spi_host0_sd_p2d,
  output logic       cio_spi_host0_sck_d2p,
  output logic       cio_spi_host0_sck_en_d2p,
  output logic       cio_spi_host0_csb_d2p,
  output logic       cio_spi_host0_csb_en_d2p,
  output logic [3:0] cio_spi_host0_sd_d2p,
  output logic [3:0] cio_spi_host0_sd_en_d2p,
  // spi_host1
  input logic [3:0]  cio_spi_host1_sd_p2d,
  output logic       cio_spi_host1_sck_d2p,
  output logic       cio_spi_host1_sck_en_d2p,
  output logic       cio_spi_host1_csb_d2p,
  output logic       cio_spi_host1_csb_en_d2p,
  output logic [3:0] cio_spi_host1_sd_d2p,
  output logic [3:0] cio_spi_host1_sd_en_d2p,

  // pad attributes to padring
  output             prim_pad_wrapper_pkg::pad_attr_t [pinmux_reg_pkg::NMioPads-1:0] mio_attr_o,
  output             prim_pad_wrapper_pkg::pad_attr_t [pinmux_reg_pkg::NDioPads-1:0] dio_attr_o,


  // Inter-module Signal External type
  output             ast_pkg::adc_ast_req_t adc_req_o,
  input              ast_pkg::adc_ast_rsp_t adc_rsp_i,
  input              edn_pkg::edn_req_t ast_edn_req_i,
  
  output             edn_pkg::edn_rsp_t ast_edn_rsp_o,
  output             lc_ctrl_pkg::lc_tx_t ast_lc_dft_en_o,
  
  input              prim_ram_1p_pkg::ram_1p_cfg_t ram_1p_cfg_i,
  input              prim_ram_2p_pkg::ram_2p_cfg_t ram_2p_cfg_i,
  input              prim_rom_pkg::rom_cfg_t rom_cfg_i,
  
  input logic        clk_main_i,
  input logic        clk_io_i,
  input logic        clk_usb_i,
  input logic        clk_aon_i,
  output logic       clk_main_jitter_en_o,
  
  output             lc_ctrl_pkg::lc_tx_t ast_clk_byp_req_o,
  input              lc_ctrl_pkg::lc_tx_t ast_clk_byp_ack_i,
  
  output             ast_pkg::ast_dif_t flash_alert_o,
  input              lc_ctrl_pkg::lc_tx_t flash_bist_enable_i,
  input logic        flash_power_down_h_i,
  input logic        flash_power_ready_h_i,
  inout [1:0]        flash_test_mode_a_io,
  inout              flash_test_voltage_h_io,
  
  output             entropy_src_pkg::entropy_src_rng_req_t es_rng_req_o,
  input              entropy_src_pkg::entropy_src_rng_rsp_t es_rng_rsp_i,
  output logic       es_rng_fips_o,
  
  output             tlul_pkg::tl_h2d_t ast_tl_req_o,
  input              tlul_pkg::tl_d2h_t ast_tl_rsp_i,
  
  output             pinmux_pkg::dft_strap_test_req_t dft_strap_test_o,
  input logic        dft_hold_tap_sel_i,
   
  output             otp_ctrl_pkg::otp_ast_req_t otp_ctrl_otp_ast_pwr_seq_o,
  input              otp_ctrl_pkg::otp_ast_rsp_t otp_ctrl_otp_ast_pwr_seq_h_i,
  inout              otp_ext_voltage_h_io,
  output             ast_pkg::ast_dif_t otp_alert_o,
  
  input logic        por_n_i,
  
  input              ast_pkg::ast_alert_req_t sensor_ctrl_ast_alert_req_i,
  output             ast_pkg::ast_alert_rsp_t sensor_ctrl_ast_alert_rsp_o,
  input              ast_pkg::ast_status_t sensor_ctrl_ast_status_i,
  input logic [8:0]  ast2pinmux_i,
  input logic        ast_init_done_i,
  
  output logic       usbdev_usb_ref_val_o,
  output logic       usbdev_usb_ref_pulse_o,
  
  output             clkmgr_pkg::clkmgr_ast_out_t clks_ast_o,
  output             rstmgr_pkg::rstmgr_ast_out_t rsts_ast_o,
  
  output logic       test_reset,
   
  output             axi_req_t axi_req,
  input              axi_resp_t axi_rsp,

  input logic        irq_ibex_i,

  input              scan_rst_ni, // reset used for test mode
  input              scan_en_i,
  input              lc_ctrl_pkg::lc_tx_t scanmode_i,   // lc_ctrl_pkg::On for Scan
   
  input              jtag_pkg::jtag_req_t jtag_i,
  output             jtag_pkg::jtag_rsp_t jtag_o,

  input logic        rst_ibex_n
  );
  
   
    
  localparam int NrDevices = 3;
  localparam int NrHosts = 1;

  import tlul_pkg::*;
  import top_pkg::*;
  import tl_main_pkg::*;
  import top_earlgrey_pkg::*;
  // Compile-time random constants
  import top_earlgrey_rnd_cnst_pkg::*;

  
  pwrmgr_pkg::pwr_ast_req_t pwrmgr_ast_req_o;
  pwrmgr_pkg::pwr_ast_rsp_t pwrmgr_ast_rsp_i = '1;

  //pwrmgr_ast_rsp_i.main_pok = 1'b1;
   
   
    
  // Test Reset to provide as output to alsaqr to start the boot
  logic trigger;
  logic [31:0] count;
  logic t_enable;
 
  enum {HIGH, LOW} state, next_state;

  always_ff @(posedge clk_main_i, negedge por_n_i) begin
		if(por_n_i == 0)
			state <= LOW;
		else
	    state <= next_state;
	end
   
  always_comb begin
	    
    trigger  = 1'b0;
    t_enable = 1'b1;
     
		case(state)
      
			LOW:      if(count == 31'b10000)
						      next_state = HIGH;
					      else 					      
                	next_state = LOW;

		  HIGH:     begin
	              trigger  = 1'b1;                
                t_enable = 1'b0;
                end
      
			default:  next_state = LOW;
      
		endcase
	end // always_comb

  assign test_reset = trigger;
  

	always_ff @(posedge clk_main_i, negedge por_n_i)
	begin
		if(por_n_i == 0)
			  count <= 'b0;
		else
			if(t_enable)
				count <= count + 1;
			else	
				count <= 'b0;
	end
 
  localparam logic [31:0] JTAG_IDCODE = {
    4'h0,     // Version
    16'h4F54, // Part Number: "OT"
    11'h426,  // Manufacturer Identity: Google
    1'b1      // (fixed)
  };

   // Signals
  logic [54:0] mio_p2d;
  logic [74:0] mio_d2p;
  logic [74:0] mio_en_d2p;
  logic [23:0] dio_p2d;
  logic [23:0] dio_d2p;
  logic [23:0] dio_en_d2p;
  // uart0
  logic        cio_uart0_rx_p2d;
  logic        cio_uart0_tx_d2p;
  logic        cio_uart0_tx_en_d2p;
  // uart1
  logic        cio_uart1_rx_p2d;
  logic        cio_uart1_tx_d2p;
  logic        cio_uart1_tx_en_d2p;
  // uart2
  logic        cio_uart2_rx_p2d;
  logic        cio_uart2_tx_d2p;
  logic        cio_uart2_tx_en_d2p;
  // uart3
  logic        cio_uart3_rx_p2d;
  logic        cio_uart3_tx_d2p;
  logic        cio_uart3_tx_en_d2p;
  // gpio
  logic [31:0] cio_gpio_gpio_p2d;
  logic [31:0] cio_gpio_gpio_d2p;
  logic [31:0] cio_gpio_gpio_en_d2p;
  
  // i2c0
  logic        cio_i2c0_sda_p2d;
  logic        cio_i2c0_scl_p2d;
  logic        cio_i2c0_sda_d2p;
  logic        cio_i2c0_sda_en_d2p;
  logic        cio_i2c0_scl_d2p;
  logic        cio_i2c0_scl_en_d2p;
  // i2c1
  logic        cio_i2c1_sda_p2d;
  logic        cio_i2c1_scl_p2d;
  logic        cio_i2c1_sda_d2p;
  logic        cio_i2c1_sda_en_d2p;
  logic        cio_i2c1_scl_d2p;
  logic        cio_i2c1_scl_en_d2p;
  // i2c2
  logic        cio_i2c2_sda_p2d;
  logic        cio_i2c2_scl_p2d;
  logic        cio_i2c2_sda_d2p;
  logic        cio_i2c2_sda_en_d2p;
  logic        cio_i2c2_scl_d2p;
  logic        cio_i2c2_scl_en_d2p;
  // pattgen
  logic        cio_pattgen_pda0_tx_d2p;
  logic        cio_pattgen_pda0_tx_en_d2p;
  logic        cio_pattgen_pcl0_tx_d2p;
  logic        cio_pattgen_pcl0_tx_en_d2p;
  logic        cio_pattgen_pda1_tx_d2p;
  logic        cio_pattgen_pda1_tx_en_d2p;
  logic        cio_pattgen_pcl1_tx_d2p;
  logic        cio_pattgen_pcl1_tx_en_d2p;
  // rv_timer
  // usbdev
  logic        cio_usbdev_sense_p2d;
  logic        cio_usbdev_d_p2d;
  logic        cio_usbdev_dp_p2d;
  logic        cio_usbdev_dn_p2d;
  logic        cio_usbdev_se0_d2p;
  logic        cio_usbdev_se0_en_d2p;
  logic        cio_usbdev_dp_pullup_d2p;
  logic        cio_usbdev_dp_pullup_en_d2p;
  logic        cio_usbdev_dn_pullup_d2p;
  logic        cio_usbdev_dn_pullup_en_d2p;
  logic        cio_usbdev_tx_mode_se_d2p;
  logic        cio_usbdev_tx_mode_se_en_d2p;
  logic        cio_usbdev_suspend_d2p;
  logic        cio_usbdev_suspend_en_d2p;
  logic        cio_usbdev_rx_enable_d2p;
  logic        cio_usbdev_rx_enable_en_d2p;
  logic        cio_usbdev_d_d2p;
  logic        cio_usbdev_d_en_d2p;
  logic        cio_usbdev_dp_d2p;
  logic        cio_usbdev_dp_en_d2p;
  logic        cio_usbdev_dn_d2p;
  logic        cio_usbdev_dn_en_d2p;
  // otp_ctrl
  logic [7:0]  cio_otp_ctrl_test_d2p;
  logic [7:0]  cio_otp_ctrl_test_en_d2p;
  // lc_ctrl
  // alerthandler
  // pwrmgr_aon
  // rstmgr_aon
  // clkmgr_aon
  // sysrst_ctrl_aon
  logic        cio_sysrst_ctrl_aon_ac_present_p2d;
  logic        cio_sysrst_ctrl_aon_key0_in_p2d;
  logic        cio_sysrst_ctrl_aon_key1_in_p2d;
  logic        cio_sysrst_ctrl_aon_key2_in_p2d;
  logic        cio_sysrst_ctrl_aon_pwrb_in_p2d;
  logic        cio_sysrst_ctrl_aon_lid_open_p2d;
  logic        cio_sysrst_ctrl_aon_ec_rst_l_p2d;
  logic        cio_sysrst_ctrl_aon_bat_disable_d2p;
  logic        cio_sysrst_ctrl_aon_bat_disable_en_d2p;
  logic        cio_sysrst_ctrl_aon_flash_wp_l_d2p;
  logic        cio_sysrst_ctrl_aon_flash_wp_l_en_d2p;
  logic        cio_sysrst_ctrl_aon_key0_out_d2p;
  logic        cio_sysrst_ctrl_aon_key0_out_en_d2p;
  logic        cio_sysrst_ctrl_aon_key1_out_d2p;
  logic        cio_sysrst_ctrl_aon_key1_out_en_d2p;
  logic        cio_sysrst_ctrl_aon_key2_out_d2p;
  logic        cio_sysrst_ctrl_aon_key2_out_en_d2p;
  logic        cio_sysrst_ctrl_aon_pwrb_out_d2p;
  logic        cio_sysrst_ctrl_aon_pwrb_out_en_d2p;
  logic        cio_sysrst_ctrl_aon_z3_wakeup_d2p;
  logic        cio_sysrst_ctrl_aon_z3_wakeup_en_d2p;
  logic        cio_sysrst_ctrl_aon_ec_rst_l_d2p;
  logic        cio_sysrst_ctrl_aon_ec_rst_l_en_d2p;
  // adc_ctrl_aon
  // pwm_aon
  logic [5:0]  cio_pwm_aon_pwm_d2p;
  logic [5:0]  cio_pwm_aon_pwm_en_d2p;
  // pinmux_aon
  // aon_timer_aon
  // sensor_ctrl_aon
  logic [8:0]  cio_sensor_ctrl_aon_ast_debug_out_d2p;
  logic [8:0]  cio_sensor_ctrl_aon_ast_debug_out_en_d2p;
  // sram_ctrl_ret_aon
  // flash_ctrl
  logic        cio_flash_ctrl_tck_p2d;
  logic        cio_flash_ctrl_tms_p2d;
  logic        cio_flash_ctrl_tdi_p2d;
  logic        cio_flash_ctrl_tdo_d2p;
  logic        cio_flash_ctrl_tdo_en_d2p;
  // rv_dm
  // rv_plic
  // aes
  // hmac
  // kmac
  // keymgr
  // csrng
  // entropy_src
  // edn0
  // edn1
  // sram_ctrl_main
  // otbn
  // rom_ctrl
  // rv_core_ibex


  logic [179:0]  intr_vector;
  // Interrupt source list
  logic intr_uart0_tx_watermark;
  logic intr_uart0_rx_watermark;
  logic intr_uart0_tx_empty;
  logic intr_uart0_rx_overflow;
  logic intr_uart0_rx_frame_err;
  logic intr_uart0_rx_break_err;
  logic intr_uart0_rx_timeout;
  logic intr_uart0_rx_parity_err;
  logic intr_uart1_tx_watermark;
  logic intr_uart1_rx_watermark;
  logic intr_uart1_tx_empty;
  logic intr_uart1_rx_overflow;
  logic intr_uart1_rx_frame_err;
  logic intr_uart1_rx_break_err;
  logic intr_uart1_rx_timeout;
  logic intr_uart1_rx_parity_err;
  logic intr_uart2_tx_watermark;
  logic intr_uart2_rx_watermark;
  logic intr_uart2_tx_empty;
  logic intr_uart2_rx_overflow;
  logic intr_uart2_rx_frame_err;
  logic intr_uart2_rx_break_err;
  logic intr_uart2_rx_timeout;
  logic intr_uart2_rx_parity_err;
  logic intr_uart3_tx_watermark;
  logic intr_uart3_rx_watermark;
  logic intr_uart3_tx_empty;
  logic intr_uart3_rx_overflow;
  logic intr_uart3_rx_frame_err;
  logic intr_uart3_rx_break_err;
  logic intr_uart3_rx_timeout;
  logic intr_uart3_rx_parity_err;
  logic [31:0] intr_gpio_gpio;
  logic intr_spi_device_rxf;
  logic intr_spi_device_rxlvl;
  logic intr_spi_device_txlvl;
  logic intr_spi_device_rxerr;
  logic intr_spi_device_rxoverflow;
  logic intr_spi_device_txunderflow;
  logic intr_spi_host0_error;
  logic intr_spi_host0_spi_event;
  logic intr_spi_host1_error;
  logic intr_spi_host1_spi_event;
  logic intr_i2c0_fmt_watermark;
  logic intr_i2c0_rx_watermark;
  logic intr_i2c0_fmt_overflow;
  logic intr_i2c0_rx_overflow;
  logic intr_i2c0_nak;
  logic intr_i2c0_scl_interference;
  logic intr_i2c0_sda_interference;
  logic intr_i2c0_stretch_timeout;
  logic intr_i2c0_sda_unstable;
  logic intr_i2c0_trans_complete;
  logic intr_i2c0_tx_empty;
  logic intr_i2c0_tx_nonempty;
  logic intr_i2c0_tx_overflow;
  logic intr_i2c0_acq_overflow;
  logic intr_i2c0_ack_stop;
  logic intr_i2c0_host_timeout;
  logic intr_i2c1_fmt_watermark;
  logic intr_i2c1_rx_watermark;
  logic intr_i2c1_fmt_overflow;
  logic intr_i2c1_rx_overflow;
  logic intr_i2c1_nak;
  logic intr_i2c1_scl_interference;
  logic intr_i2c1_sda_interference;
  logic intr_i2c1_stretch_timeout;
  logic intr_i2c1_sda_unstable;
  logic intr_i2c1_trans_complete;
  logic intr_i2c1_tx_empty;
  logic intr_i2c1_tx_nonempty;
  logic intr_i2c1_tx_overflow;
  logic intr_i2c1_acq_overflow;
  logic intr_i2c1_ack_stop;
  logic intr_i2c1_host_timeout;
  logic intr_i2c2_fmt_watermark;
  logic intr_i2c2_rx_watermark;
  logic intr_i2c2_fmt_overflow;
  logic intr_i2c2_rx_overflow;
  logic intr_i2c2_nak;
  logic intr_i2c2_scl_interference;
  logic intr_i2c2_sda_interference;
  logic intr_i2c2_stretch_timeout;
  logic intr_i2c2_sda_unstable;
  logic intr_i2c2_trans_complete;
  logic intr_i2c2_tx_empty;
  logic intr_i2c2_tx_nonempty;
  logic intr_i2c2_tx_overflow;
  logic intr_i2c2_acq_overflow;
  logic intr_i2c2_ack_stop;
  logic intr_i2c2_host_timeout;
  logic intr_pattgen_done_ch0;
  logic intr_pattgen_done_ch1;
  logic intr_rv_timer_timer_expired_0_0;
  logic intr_usbdev_pkt_received;
  logic intr_usbdev_pkt_sent;
  logic intr_usbdev_disconnected;
  logic intr_usbdev_host_lost;
  logic intr_usbdev_link_reset;
  logic intr_usbdev_link_suspend;
  logic intr_usbdev_link_resume;
  logic intr_usbdev_av_empty;
  logic intr_usbdev_rx_full;
  logic intr_usbdev_av_overflow;
  logic intr_usbdev_link_in_err;
  logic intr_usbdev_rx_crc_err;
  logic intr_usbdev_rx_pid_err;
  logic intr_usbdev_rx_bitstuff_err;
  logic intr_usbdev_frame;
  logic intr_usbdev_connected;
  logic intr_usbdev_link_out_err;
  logic intr_otp_ctrl_otp_operation_done;
  logic intr_otp_ctrl_otp_error;
  logic intr_alert_handler_classa;
  logic intr_alert_handler_classb;
  logic intr_alert_handler_classc;
  logic intr_alert_handler_classd;
  logic intr_pwrmgr_aon_wakeup;
  logic intr_sysrst_ctrl_aon_sysrst_ctrl;
  logic intr_adc_ctrl_aon_debug_cable;
  logic intr_aon_timer_aon_wkup_timer_expired;
  logic intr_aon_timer_aon_wdog_timer_bark;
  logic intr_flash_ctrl_prog_empty;
  logic intr_flash_ctrl_prog_lvl;
  logic intr_flash_ctrl_rd_full;
  logic intr_flash_ctrl_rd_lvl;
  logic intr_flash_ctrl_op_done;
  logic intr_flash_ctrl_err;
  logic intr_hmac_hmac_done;
  logic intr_hmac_fifo_empty;
  logic intr_hmac_hmac_err;
  logic intr_kmac_kmac_done;
  logic intr_kmac_fifo_empty;
  logic intr_kmac_kmac_err;
  logic intr_keymgr_op_done;
  logic intr_csrng_cs_cmd_req_done;
  logic intr_csrng_cs_entropy_req;
  logic intr_csrng_cs_hw_inst_exc;
  logic intr_csrng_cs_fatal_err;
  logic intr_entropy_src_es_entropy_valid;
  logic intr_entropy_src_es_health_test_failed;
  logic intr_entropy_src_es_observe_fifo_ready;
  logic intr_entropy_src_es_fatal_err;
  logic intr_edn0_edn_cmd_req_done;
  logic intr_edn0_edn_fatal_err;
  logic intr_edn1_edn_cmd_req_done;
  logic intr_edn1_edn_fatal_err;
  logic intr_otbn_done;

  // simctrl signals
  logic           device_req;
  logic [31:0]    device_addr;
  logic           device_we;
  logic [ 3:0]    device_be;
  logic [31:0]    device_wdata;
  logic           device_rvalid; 
  logic [31:0]    device_rdata;
  logic           device_err;

  // simcontrol ibexprot2tlul
   
   assign device_req             = core2simctrl.a_valid;
   assign device_addr            = core2simctrl.a_address;
   assign device_be              = core2simctrl.a_mask;
   assign device_we              =  ~(core2simctrl.a_opcode[2] || core2simctrl.a_opcode[0]);
   assign device_wdata           = core2simctrl.a_data;
   assign simctrl2core.d_valid   = device_rvalid; 
   assign simctrl2core.a_ready   = 1'b1; 
   assign simctrl2core.d_data    = device_rdata;
   assign simctrl2core.d_opcode  = tlul_pkg::AccessAckData;
   assign simctrl2core.d_error   = device_err;
   assign simctrl2core.d_param   = core2simctrl.a_param;
   assign simctrl2core.d_size    = core2simctrl.a_size;
   assign simctrl2core.d_source  = core2simctrl.a_source;
   assign simctrl2core.d_user    = TL_D_USER_DEFAULT;
   assign simctrl2core.d_sink    = '0;

   assign device_err = 1'b0;

  

/*     
  typedef enum logic[1:0] {
    Ram,
    SimCtrl,
    Timer
  } bus_device_e;

  // host and device signals
  logic           host_req    [NrHosts]; 
  logic           host_gnt    [NrHosts];
  logic [31:0]    host_addr   [NrHosts]; 
  logic           host_we     [NrHosts];
  logic [ 3:0]    host_be     [NrHosts];
  logic [31:0]    host_wdata  [NrHosts];
  logic           host_rvalid [NrHosts];
  logic [31:0]    host_rdata  [NrHosts];
  logic           host_err    [NrHosts];

  // devices (slaves)
  logic           device_req    [NrDevices];
  logic [31:0]    device_addr   [NrDevices];
  logic           device_we     [NrDevices];
  logic [ 3:0]    device_be     [NrDevices];
  logic [31:0]    device_wdata  [NrDevices];
  logic           device_rvalid [NrDevices]; 
  logic [31:0]    device_rdata  [NrDevices];
  logic           device_err    [NrDevices];

  logic           device_req_;
  logic [31:0]    device_addr_;
  logic           device_we_;
  logic [ 3:0]    device_be_;
  logic [31:0]    device_wdata_;
  logic           device_rvalid_; 
  logic [31:0]    device_rdata_;
  logic           device_err_;
   

  // Instruction fetch signals
  logic instr_req;
  logic instr_gnt;
  logic instr_rvalid;
  logic [31:0] instr_addr;
  logic [31:0] instr_rdata;
  logic instr_err;

  assign instr_gnt = instr_req;
  assign instr_err = '0;

 

  // Tie-off unused error signals
  assign device_err[Ram] = 1'b0;
  assign device_err_     = 1'b0;
  assign device_err[SimCtrl] = 1'b0;

// protocol conversion for the simctrl and ram, not opentitan ips so not implementing tile link
// instructions interface

    tlul_pkg::tl_d_user_t                  tieoff;
   
    assign instr_req                       = core2instr.a_valid;
    assign instr_addr                      = core2instr.a_address;
    assign instr2core.d_valid              = instr_rvalid; 
    assign instr2core.d_data               = instr_rdata;
    assign instr2core.a_ready              = 1'b1;
    assign instr2core.d_error              = instr_err;
    assign instr2core.d_opcode             = tlul_pkg::AccessAckData;  
    assign instr2core.d_param              = core2instr.a_param;
    assign instr2core.d_size               = core2instr.a_size;
    assign instr2core.d_source             = core2instr.a_source;
    assign instr2core.d_sink               = '0;
    assign instr2core.d_user               = TL_D_USER_DEFAULT;
 


  
// simcontrol ibexprot2tlul
   
    assign device_req[SimCtrl]             = core2simctrl.a_valid;
    assign device_addr[SimCtrl]            = core2simctrl.a_address;
    assign device_be[SimCtrl]              = core2simctrl.a_mask;
    assign device_we[SimCtrl]              =  ~(core2simctrl.a_opcode[2] || core2simctrl.a_opcode[0]);
    assign device_wdata[SimCtrl]           = core2simctrl.a_data;
    assign simctrl2core.d_valid            = device_rvalid[SimCtrl]; 
    assign simctrl2core.a_ready            = 1'b1; 
    assign simctrl2core.d_data             = device_rdata[SimCtrl];
    assign simctrl2core.d_opcode           = tlul_pkg::AccessAckData;
    assign simctrl2core.d_error            = device_err[SimCtrl];
    assign simctrl2core.d_param            = core2simctrl.a_param;
    assign simctrl2core.d_size             = core2simctrl.a_size;
    assign simctrl2core.d_source           = core2simctrl.a_source;
    assign simctrl2core.d_user             = TL_D_USER_DEFAULT;
    assign simctrl2core.d_sink               = '0;

// test ram ibexprot2tlul
   
    assign device_req_              = tcore2simctrl.a_valid;
    assign device_addr_             = tcore2simctrl.a_address;
    assign device_be_               = tcore2simctrl.a_mask;
    assign device_we_               =  ~(tcore2simctrl.a_opcode[2] || tcore2simctrl.a_opcode[0]);
    assign device_wdata_            = tcore2simctrl.a_data;
    assign tsimctrl2core.d_valid    = device_rvalid_; 
    assign tsimctrl2core.a_ready    = 1'b1; 
    assign tsimctrl2core.d_data     = device_rdata_;
    assign tsimctrl2core.d_opcode   = tlul_pkg::AccessAckData;
    assign tsimctrl2core.d_error    = device_err_;
    assign tsimctrl2core.d_param    = tcore2simctrl.a_param;
    assign tsimctrl2core.d_size     = tcore2simctrl.a_size;
    assign tsimctrl2core.d_source   = tcore2simctrl.a_source;
    assign tsimctrl2core.d_user     = TL_D_USER_DEFAULT;
    assign tsimctrl2core.d_sink     = '0; 


// ram ibexprot2tlul
   
    assign device_req[Ram]                 = core2ram.a_valid;
    assign device_addr[Ram]                = core2ram.a_address;
    assign device_be[Ram]                  = core2ram.a_mask;
    assign device_we[Ram]                  =  ~(core2ram.a_opcode[2] ||  core2ram.a_opcode[0]);
    assign device_wdata[Ram]               = core2ram.a_data;
    assign ram2core.d_valid                = device_rvalid[Ram]; 
    assign ram2core.a_ready                = 1'b1; 
    assign ram2core.d_data                 = device_rdata[Ram];
    assign ram2core.d_opcode               = tlul_pkg::AccessAckData;
    assign ram2core.d_error                = device_err[Ram];
    assign ram2core.d_param                = core2ram.a_param;
    assign ram2core.d_size                 = core2ram.a_size;
    assign ram2core.d_source               = core2ram.a_source;
    assign ram2core.d_user                 = TL_D_USER_DEFAULT;
    assign ram2core.d_sink                 = '0;
   
*/   
  // Alert list
  prim_alert_pkg::alert_tx_t [alert_pkg::NAlerts-1:0]  alert_tx;
  prim_alert_pkg::alert_rx_t [alert_pkg::NAlerts-1:0]  alert_rx;


  // define inter-module signals
  prim_ram_1p_pkg::ram_1p_cfg_t       ast_ram_1p_cfg;
  prim_ram_2p_pkg::ram_2p_cfg_t       ast_ram_2p_cfg;
  prim_rom_pkg::rom_cfg_t       ast_rom_cfg;
  alert_pkg::alert_crashdump_t       alert_handler_crashdump;
  prim_esc_pkg::esc_rx_t [3:0] alert_handler_esc_rx;
  prim_esc_pkg::esc_tx_t [3:0] alert_handler_esc_tx;
  logic       aon_timer_aon_nmi_wdog_timer_bark;
  csrng_pkg::csrng_req_t [1:0] csrng_csrng_cmd_req;
  csrng_pkg::csrng_rsp_t [1:0] csrng_csrng_cmd_rsp;
  entropy_src_pkg::entropy_src_hw_if_req_t       csrng_entropy_src_hw_if_req;
  entropy_src_pkg::entropy_src_hw_if_rsp_t       csrng_entropy_src_hw_if_rsp;
  entropy_src_pkg::cs_aes_halt_req_t       csrng_cs_aes_halt_req;
  entropy_src_pkg::cs_aes_halt_rsp_t       csrng_cs_aes_halt_rsp;
  flash_ctrl_pkg::keymgr_flash_t       flash_ctrl_keymgr;
  otp_ctrl_pkg::flash_otp_key_req_t       flash_ctrl_otp_req;
  otp_ctrl_pkg::flash_otp_key_rsp_t       flash_ctrl_otp_rsp;
  lc_ctrl_pkg::lc_tx_t       flash_ctrl_rma_req;
  lc_ctrl_pkg::lc_tx_t       flash_ctrl_rma_ack;
  lc_ctrl_pkg::lc_flash_rma_seed_t       flash_ctrl_rma_seed;
  otp_ctrl_pkg::sram_otp_key_req_t [1:0] otp_ctrl_sram_otp_key_req;
  otp_ctrl_pkg::sram_otp_key_rsp_t [1:0] otp_ctrl_sram_otp_key_rsp;
  pwrmgr_pkg::pwr_flash_t       pwrmgr_aon_pwr_flash;
  pwrmgr_pkg::pwr_rst_req_t       pwrmgr_aon_pwr_rst_req;
  pwrmgr_pkg::pwr_rst_rsp_t       pwrmgr_aon_pwr_rst_rsp;
  pwrmgr_pkg::pwr_clk_req_t       pwrmgr_aon_pwr_clk_req;
  pwrmgr_pkg::pwr_clk_rsp_t       pwrmgr_aon_pwr_clk_rsp;
  pwrmgr_pkg::pwr_otp_req_t       pwrmgr_aon_pwr_otp_req;
  pwrmgr_pkg::pwr_otp_rsp_t       pwrmgr_aon_pwr_otp_rsp;
  pwrmgr_pkg::pwr_lc_req_t       pwrmgr_aon_pwr_lc_req;
  pwrmgr_pkg::pwr_lc_rsp_t       pwrmgr_aon_pwr_lc_rsp;
  logic       pwrmgr_aon_strap;
  logic       pwrmgr_aon_low_power;
  lc_ctrl_pkg::lc_tx_t       pwrmgr_aon_fetch_en;
  rom_ctrl_pkg::pwrmgr_data_t       rom_ctrl_pwrmgr_data;
  rom_ctrl_pkg::keymgr_data_t       rom_ctrl_keymgr_data;
  logic       usbdev_usb_out_of_rst;
  logic       usbdev_usb_aon_wake_en;
  logic       usbdev_usb_aon_wake_ack;
  logic       usbdev_usb_suspend;
  usbdev_pkg::awk_state_t       pinmux_aon_usb_state_debug;
  edn_pkg::edn_req_t [6:0] edn0_edn_req;
  edn_pkg::edn_rsp_t [6:0] edn0_edn_rsp;
  edn_pkg::edn_req_t [6:0] edn1_edn_req;
  edn_pkg::edn_rsp_t [6:0] edn1_edn_rsp;
  otp_ctrl_pkg::otbn_otp_key_req_t       otp_ctrl_otbn_otp_key_req;
  otp_ctrl_pkg::otbn_otp_key_rsp_t       otp_ctrl_otbn_otp_key_rsp;
  otp_ctrl_pkg::otp_keymgr_key_t       otp_ctrl_otp_keymgr_key;
  keymgr_pkg::hw_key_req_t       keymgr_kmac_key;
  kmac_pkg::app_req_t [2:0] kmac_app_req;
  kmac_pkg::app_rsp_t [2:0] kmac_app_rsp;
  logic       kmac_en_masking;
  logic [4:0] clkmgr_aon_idle;
  jtag_pkg::jtag_req_t       pinmux_aon_lc_jtag_req;
  jtag_pkg::jtag_rsp_t       pinmux_aon_lc_jtag_rsp;
  jtag_pkg::jtag_req_t       pinmux_aon_rv_jtag_req;
  jtag_pkg::jtag_rsp_t       pinmux_aon_rv_jtag_rsp;
  otp_ctrl_pkg::otp_lc_data_t       otp_ctrl_otp_lc_data;
  otp_ctrl_pkg::lc_otp_program_req_t       lc_ctrl_lc_otp_program_req;
  otp_ctrl_pkg::lc_otp_program_rsp_t       lc_ctrl_lc_otp_program_rsp;
  otp_ctrl_pkg::lc_otp_vendor_test_req_t       lc_ctrl_lc_otp_vendor_test_req;
  otp_ctrl_pkg::lc_otp_vendor_test_rsp_t       lc_ctrl_lc_otp_vendor_test_rsp;
  lc_ctrl_pkg::lc_keymgr_div_t       lc_ctrl_lc_keymgr_div;
  lc_ctrl_pkg::lc_tx_t       lc_ctrl_lc_dft_en;
  lc_ctrl_pkg::lc_tx_t       lc_ctrl_lc_nvm_debug_en;
  lc_ctrl_pkg::lc_tx_t       lc_ctrl_lc_hw_debug_en;
  lc_ctrl_pkg::lc_tx_t       lc_ctrl_lc_cpu_en;
  lc_ctrl_pkg::lc_tx_t       lc_ctrl_lc_keymgr_en;
  lc_ctrl_pkg::lc_tx_t       lc_ctrl_lc_escalate_en;
  lc_ctrl_pkg::lc_tx_t       lc_ctrl_lc_check_byp_en;
  lc_ctrl_pkg::lc_tx_t       lc_ctrl_lc_clk_byp_req;
  lc_ctrl_pkg::lc_tx_t       lc_ctrl_lc_clk_byp_ack;
  lc_ctrl_pkg::lc_tx_t       lc_ctrl_lc_creator_seed_sw_rw_en;
  lc_ctrl_pkg::lc_tx_t       lc_ctrl_lc_owner_seed_sw_rw_en;
  lc_ctrl_pkg::lc_tx_t       lc_ctrl_lc_iso_part_sw_rd_en;
  lc_ctrl_pkg::lc_tx_t       lc_ctrl_lc_iso_part_sw_wr_en;
  lc_ctrl_pkg::lc_tx_t       lc_ctrl_lc_seed_hw_rd_en;
  logic       rv_plic_msip;
  logic       rv_plic_irq;
  logic       rv_dm_debug_req;
  logic       rv_core_ibex_rst_cpu_n;
  ibex_pkg::crash_dump_t       rv_core_ibex_crash_dump;
  pwrmgr_pkg::pwr_cpu_t       rv_core_ibex_pwrmgr;
  spi_device_pkg::passthrough_req_t       spi_device_passthrough_req;
  spi_device_pkg::passthrough_rsp_t       spi_device_passthrough_rsp;
  logic       rv_dm_ndmreset_req;
  logic [4:0] pwrmgr_aon_wakeups;
  logic [1:0] pwrmgr_aon_rstreqs;

   
  tlul_pkg::tl_h2d_t       main_tl_rv_core_ibex__corei_req;
  tlul_pkg::tl_d2h_t       main_tl_rv_core_ibex__corei_rsp;
  tlul_pkg::tl_h2d_t       main_tl_rv_core_ibex__cored_req;
  tlul_pkg::tl_d2h_t       main_tl_rv_core_ibex__cored_rsp;
  tlul_pkg::tl_h2d_t       main_tl_rv_dm__sba_req;
  tlul_pkg::tl_d2h_t       main_tl_rv_dm__sba_rsp;
  tlul_pkg::tl_h2d_t       rv_dm_regs_tl_d_req;
  tlul_pkg::tl_d2h_t       rv_dm_regs_tl_d_rsp;
  tlul_pkg::tl_h2d_t       rv_dm_rom_tl_d_req;
  tlul_pkg::tl_d2h_t       rv_dm_rom_tl_d_rsp;
  tlul_pkg::tl_h2d_t       rom_ctrl_rom_tl_req;
  tlul_pkg::tl_d2h_t       rom_ctrl_rom_tl_rsp;
  tlul_pkg::tl_h2d_t       rom_ctrl_regs_tl_req;
  tlul_pkg::tl_d2h_t       rom_ctrl_regs_tl_rsp;
  tlul_pkg::tl_h2d_t       main_tl_peri_req;
  tlul_pkg::tl_d2h_t       main_tl_peri_rsp;
  tlul_pkg::tl_h2d_t       flash_ctrl_core_tl_req;
  tlul_pkg::tl_d2h_t       flash_ctrl_core_tl_rsp;
  tlul_pkg::tl_h2d_t       flash_ctrl_prim_tl_req;
  tlul_pkg::tl_d2h_t       flash_ctrl_prim_tl_rsp;
  tlul_pkg::tl_h2d_t       flash_ctrl_mem_tl_req;
  tlul_pkg::tl_d2h_t       flash_ctrl_mem_tl_rsp;
  tlul_pkg::tl_h2d_t       hmac_tl_req;
  tlul_pkg::tl_d2h_t       hmac_tl_rsp;
  tlul_pkg::tl_h2d_t       kmac_tl_req;
  tlul_pkg::tl_d2h_t       kmac_tl_rsp;
  tlul_pkg::tl_h2d_t       aes_tl_req;
  tlul_pkg::tl_d2h_t       aes_tl_rsp;
  tlul_pkg::tl_h2d_t       entropy_src_tl_req;
  tlul_pkg::tl_d2h_t       entropy_src_tl_rsp;
  tlul_pkg::tl_h2d_t       csrng_tl_req;
  tlul_pkg::tl_d2h_t       csrng_tl_rsp;
  tlul_pkg::tl_h2d_t       edn0_tl_req;
  tlul_pkg::tl_d2h_t       edn0_tl_rsp;
  tlul_pkg::tl_h2d_t       edn1_tl_req;
  tlul_pkg::tl_d2h_t       edn1_tl_rsp;
  tlul_pkg::tl_h2d_t       rv_plic_tl_req;
  tlul_pkg::tl_d2h_t       rv_plic_tl_rsp;
  tlul_pkg::tl_h2d_t       otbn_tl_req;
  tlul_pkg::tl_d2h_t       otbn_tl_rsp;
  tlul_pkg::tl_h2d_t       keymgr_tl_req;
  tlul_pkg::tl_d2h_t       keymgr_tl_rsp;
  tlul_pkg::tl_h2d_t       rv_core_ibex_cfg_tl_d_req;
  tlul_pkg::tl_d2h_t       rv_core_ibex_cfg_tl_d_rsp;
  tlul_pkg::tl_h2d_t       sram_ctrl_main_regs_tl_req;
  tlul_pkg::tl_d2h_t       sram_ctrl_main_regs_tl_rsp;
  tlul_pkg::tl_h2d_t       sram_ctrl_main_ram_tl_req;
  tlul_pkg::tl_d2h_t       sram_ctrl_main_ram_tl_rsp;
  tlul_pkg::tl_h2d_t       uart0_tl_req;
  tlul_pkg::tl_d2h_t       uart0_tl_rsp;
  tlul_pkg::tl_h2d_t       uart1_tl_req;
  tlul_pkg::tl_d2h_t       uart1_tl_rsp;
  tlul_pkg::tl_h2d_t       uart2_tl_req;
  tlul_pkg::tl_d2h_t       uart2_tl_rsp;
  tlul_pkg::tl_h2d_t       uart3_tl_req;
  tlul_pkg::tl_d2h_t       uart3_tl_rsp;
  tlul_pkg::tl_h2d_t       i2c0_tl_req;
  tlul_pkg::tl_d2h_t       i2c0_tl_rsp;
  tlul_pkg::tl_h2d_t       i2c1_tl_req;
  tlul_pkg::tl_d2h_t       i2c1_tl_rsp;
  tlul_pkg::tl_h2d_t       i2c2_tl_req;
  tlul_pkg::tl_d2h_t       i2c2_tl_rsp;
  tlul_pkg::tl_h2d_t       pattgen_tl_req;
  tlul_pkg::tl_d2h_t       pattgen_tl_rsp;
  tlul_pkg::tl_h2d_t       pwm_aon_tl_req;
  tlul_pkg::tl_d2h_t       pwm_aon_tl_rsp;
  tlul_pkg::tl_h2d_t       gpio_tl_req;
  tlul_pkg::tl_d2h_t       gpio_tl_rsp;
  tlul_pkg::tl_h2d_t       spi_device_tl_req;
  tlul_pkg::tl_d2h_t       spi_device_tl_rsp;
  tlul_pkg::tl_h2d_t       spi_host0_tl_req;
  tlul_pkg::tl_d2h_t       spi_host0_tl_rsp;
  tlul_pkg::tl_h2d_t       spi_host1_tl_req;
  tlul_pkg::tl_d2h_t       spi_host1_tl_rsp;
  tlul_pkg::tl_h2d_t       rv_timer_tl_req;
  tlul_pkg::tl_d2h_t       rv_timer_tl_rsp;
  tlul_pkg::tl_h2d_t       usbdev_tl_req;
  tlul_pkg::tl_d2h_t       usbdev_tl_rsp;
  tlul_pkg::tl_h2d_t       pwrmgr_aon_tl_req;
  tlul_pkg::tl_d2h_t       pwrmgr_aon_tl_rsp;
  tlul_pkg::tl_h2d_t       rstmgr_aon_tl_req;
  tlul_pkg::tl_d2h_t       rstmgr_aon_tl_rsp;
  tlul_pkg::tl_h2d_t       clkmgr_aon_tl_req;
  tlul_pkg::tl_d2h_t       clkmgr_aon_tl_rsp;
  tlul_pkg::tl_h2d_t       pinmux_aon_tl_req;
  tlul_pkg::tl_d2h_t       pinmux_aon_tl_rsp;
  tlul_pkg::tl_h2d_t       otp_ctrl_core_tl_req;
  tlul_pkg::tl_d2h_t       otp_ctrl_core_tl_rsp;
  tlul_pkg::tl_h2d_t       otp_ctrl_prim_tl_req;
  tlul_pkg::tl_d2h_t       otp_ctrl_prim_tl_rsp;
  tlul_pkg::tl_h2d_t       lc_ctrl_tl_req;
  tlul_pkg::tl_d2h_t       lc_ctrl_tl_rsp;
  tlul_pkg::tl_h2d_t       sensor_ctrl_aon_tl_req;
  tlul_pkg::tl_d2h_t       sensor_ctrl_aon_tl_rsp;
  tlul_pkg::tl_h2d_t       alert_handler_tl_req;
  tlul_pkg::tl_d2h_t       alert_handler_tl_rsp;
  tlul_pkg::tl_h2d_t       sram_ctrl_ret_aon_regs_tl_req;
  tlul_pkg::tl_d2h_t       sram_ctrl_ret_aon_regs_tl_rsp;
  tlul_pkg::tl_h2d_t       sram_ctrl_ret_aon_ram_tl_req;
  tlul_pkg::tl_d2h_t       sram_ctrl_ret_aon_ram_tl_rsp;
  tlul_pkg::tl_h2d_t       aon_timer_aon_tl_req;
  tlul_pkg::tl_d2h_t       aon_timer_aon_tl_rsp;
  tlul_pkg::tl_h2d_t       sysrst_ctrl_aon_tl_req;
  tlul_pkg::tl_d2h_t       sysrst_ctrl_aon_tl_rsp;
  tlul_pkg::tl_h2d_t       adc_ctrl_aon_tl_req;
  tlul_pkg::tl_d2h_t       adc_ctrl_aon_tl_rsp;


  tlul_pkg::tl_h2d_t       core2simctrl;
  tlul_pkg::tl_d2h_t       simctrl2core;
  //tlul_pkg::tl_h2d_t       core2ram;
  //tlul_pkg::tl_d2h_t       ram2core;
  //tlul_pkg::tl_h2d_t       core2instr;
  //tlul_pkg::tl_d2h_t       instr2core;
  tlul_pkg::tl_h2d_t       core2alsaqr;
  tlul_pkg::tl_d2h_t       alsaqr2core;
  
  rstmgr_pkg::rstmgr_out_t       rstmgr_aon_resets;
  clkmgr_pkg::clkmgr_out_t       clkmgr_aon_clocks;
  logic       rv_core_ibex_irq_timer;
  logic [31:0] rv_core_ibex_hart_id;
  logic [31:0] rv_core_ibex_boot_addr;
  jtag_pkg::jtag_req_t       pinmux_aon_dft_jtag_req;
  jtag_pkg::jtag_rsp_t       pinmux_aon_dft_jtag_rsp;
  otp_ctrl_part_pkg::otp_hw_cfg_t       otp_ctrl_otp_hw_cfg;
  otp_ctrl_pkg::otp_en_t       csrng_otp_en_csrng_sw_app_read;
  otp_ctrl_pkg::otp_en_t       entropy_src_otp_en_entropy_src_fw_read;
  otp_ctrl_pkg::otp_en_t       entropy_src_otp_en_entropy_src_fw_over;
  otp_ctrl_pkg::otp_device_id_t       lc_ctrl_otp_device_id;
  otp_ctrl_pkg::otp_manuf_state_t       lc_ctrl_otp_manuf_state;
  otp_ctrl_pkg::otp_device_id_t       keymgr_otp_device_id;
  otp_ctrl_pkg::otp_en_t       sram_ctrl_main_otp_en_sram_ifetch;

  edn_pkg::edn_req_t ast_tieoff;
 
  // define mixed connection to port
  assign edn0_edn_req[2] = 1'b0;//ast_edn_req_i;
  assign ast_edn_rsp_o = edn0_edn_rsp[2];
  assign ast_lc_dft_en_o = lc_ctrl_lc_dft_en;
  assign ast_ram_1p_cfg = ram_1p_cfg_i;
  assign ast_ram_2p_cfg = ram_2p_cfg_i;
  assign ast_rom_cfg = rom_cfg_i;

  // define partial inter-module tie-off
  edn_pkg::edn_rsp_t unused_edn1_edn_rsp1;
  edn_pkg::edn_rsp_t unused_edn1_edn_rsp2;
  edn_pkg::edn_rsp_t unused_edn1_edn_rsp3;
  edn_pkg::edn_rsp_t unused_edn1_edn_rsp4;
  edn_pkg::edn_rsp_t unused_edn1_edn_rsp5;
  edn_pkg::edn_rsp_t unused_edn1_edn_rsp6;

  // assign partial inter-module tie-off
  assign unused_edn1_edn_rsp1 = edn1_edn_rsp[1];
  assign unused_edn1_edn_rsp2 = edn1_edn_rsp[2];
  assign unused_edn1_edn_rsp3 = edn1_edn_rsp[3];
  assign unused_edn1_edn_rsp4 = edn1_edn_rsp[4];
  assign unused_edn1_edn_rsp5 = edn1_edn_rsp[5];
  assign unused_edn1_edn_rsp6 = edn1_edn_rsp[6];
  assign edn1_edn_req[1] = '0;
  assign edn1_edn_req[2] = '0;
  assign edn1_edn_req[3] = '0;
  assign edn1_edn_req[4] = '0;
  assign edn1_edn_req[5] = '0;
  assign edn1_edn_req[6] = '0;

  // OTP HW_CFG Broadcast signals.
  // TODO(#6713): The actual struct breakout and mapping currently needs to
  // be performed by hand.
  assign csrng_otp_en_csrng_sw_app_read = otp_ctrl_otp_hw_cfg.data.en_csrng_sw_app_read;
  assign entropy_src_otp_en_entropy_src_fw_read = otp_ctrl_otp_hw_cfg.data.en_entropy_src_fw_read;
  assign entropy_src_otp_en_entropy_src_fw_over = otp_ctrl_otp_hw_cfg.data.en_entropy_src_fw_over;
  assign sram_ctrl_main_otp_en_sram_ifetch = otp_ctrl_otp_hw_cfg.data.en_sram_ifetch;
  assign lc_ctrl_otp_device_id = otp_ctrl_otp_hw_cfg.data.device_id;
  assign lc_ctrl_otp_manuf_state = otp_ctrl_otp_hw_cfg.data.manuf_state;
  assign keymgr_otp_device_id = otp_ctrl_otp_hw_cfg.data.device_id;

  logic unused_otp_hw_cfg_bits;
  assign unused_otp_hw_cfg_bits = ^{
    otp_ctrl_otp_hw_cfg.valid,
    otp_ctrl_otp_hw_cfg.data.hw_cfg_digest,
    otp_ctrl_otp_hw_cfg.data.unallocated
  };
   
   // certain resets are unused
  logic unused_d0_rst_por_aon;
  logic unused_d0_rst_por;
  logic unused_d0_rst_por_io;
  logic unused_d0_rst_por_io_div2;
  logic unused_d0_rst_por_io_div4;
  logic unused_d0_rst_por_usb;
  logic unused_daon_rst_lc;
  logic unused_d0_rst_lc_aon;
  logic unused_daon_rst_sys;
  logic unused_daon_rst_sys_shadowed;
  logic unused_daon_rst_spi_device;
  logic unused_daon_rst_spi_host0;
  logic unused_daon_rst_spi_host0_core;
  logic unused_daon_rst_spi_host1;
  logic unused_daon_rst_spi_host1_core;
  logic unused_daon_rst_usb;
  logic unused_daon_rst_usbif;
  logic unused_daon_rst_i2c0;
  logic unused_daon_rst_i2c1;
  logic unused_daon_rst_i2c2;
  assign unused_d0_rst_por_aon = rstmgr_aon_resets.rst_por_aon_n[rstmgr_pkg::Domain0Sel];
  assign unused_d0_rst_por = rstmgr_aon_resets.rst_por_n[rstmgr_pkg::Domain0Sel];
  assign unused_d0_rst_por_io = rstmgr_aon_resets.rst_por_io_n[rstmgr_pkg::Domain0Sel];
  assign unused_d0_rst_por_io_div2 = rstmgr_aon_resets.rst_por_io_div2_n[rstmgr_pkg::Domain0Sel];
  assign unused_d0_rst_por_io_div4 = rstmgr_aon_resets.rst_por_io_div4_n[rstmgr_pkg::Domain0Sel];
  assign unused_d0_rst_por_usb = rstmgr_aon_resets.rst_por_usb_n[rstmgr_pkg::Domain0Sel];
  assign unused_daon_rst_lc = rstmgr_aon_resets.rst_lc_n[rstmgr_pkg::DomainAonSel];
  assign unused_d0_rst_lc_aon = rstmgr_aon_resets.rst_lc_aon_n[rstmgr_pkg::Domain0Sel];
  assign unused_daon_rst_sys = rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::DomainAonSel];
  assign unused_daon_rst_sys_shadowed = rstmgr_aon_resets.rst_sys_shadowed_n[rstmgr_pkg::DomainAonSel];
  assign unused_daon_rst_spi_device = rstmgr_aon_resets.rst_spi_device_n[rstmgr_pkg::DomainAonSel];
  assign unused_daon_rst_spi_host0 = rstmgr_aon_resets.rst_spi_host0_n[rstmgr_pkg::DomainAonSel];
  assign unused_daon_rst_spi_host0_core = rstmgr_aon_resets.rst_spi_host0_core_n[rstmgr_pkg::DomainAonSel];
  assign unused_daon_rst_spi_host1 = rstmgr_aon_resets.rst_spi_host1_n[rstmgr_pkg::DomainAonSel];
  assign unused_daon_rst_spi_host1_core = rstmgr_aon_resets.rst_spi_host1_core_n[rstmgr_pkg::DomainAonSel];
  assign unused_daon_rst_usb = rstmgr_aon_resets.rst_usb_n[rstmgr_pkg::DomainAonSel];
  assign unused_daon_rst_usbif = rstmgr_aon_resets.rst_usbif_n[rstmgr_pkg::DomainAonSel];
  assign unused_daon_rst_i2c0 = rstmgr_aon_resets.rst_i2c0_n[rstmgr_pkg::DomainAonSel];
  assign unused_daon_rst_i2c1 = rstmgr_aon_resets.rst_i2c1_n[rstmgr_pkg::DomainAonSel];
  assign unused_daon_rst_i2c2 = rstmgr_aon_resets.rst_i2c2_n[rstmgr_pkg::DomainAonSel];

  // ibex specific assignments
  // TODO: This should be further automated in the future.
  assign rv_core_ibex_irq_timer = intr_rv_timer_timer_expired_0_0;
  assign rv_core_ibex_hart_id = '0;
   
  assign rv_core_ibex_boot_addr = ADDR_SPACE_ROM_CTRL__ROM;

  parameter int unsigned AXI_ID_WIDTH            = 8; 
  parameter int unsigned AXI_ADDR_WIDTH          = 64; 
  parameter int unsigned AXI_SLV_PORT_DATA_WIDTH = 32; 
  parameter int unsigned AXI_MST_PORT_DATA_WIDTH = 64; 
  parameter int unsigned AXI_USER_WIDTH          = 1; 
  parameter int unsigned AXI_MAX_READS           = 1; 
 
  typedef logic [AXI_ADDR_WIDTH-1:0]            addr_t;
  typedef logic [AXI_MST_PORT_DATA_WIDTH-1:0]   data_t;
  typedef logic [AXI_MST_PORT_DATA_WIDTH/8-1:0] strb_t;

  typedef logic [AXI_ID_WIDTH-1:0] id_t                   ;
  typedef logic [AXI_MST_PORT_DATA_WIDTH-1:0] mst_data_t  ;
  typedef logic [AXI_MST_PORT_DATA_WIDTH/8-1:0] mst_strb_t;
  typedef logic [AXI_SLV_PORT_DATA_WIDTH-1:0] slv_data_t  ;
  typedef logic [AXI_SLV_PORT_DATA_WIDTH/8-1:0] slv_strb_t;
  typedef logic [AXI_USER_WIDTH-1:0] user_t;
     
  `AXI_TYPEDEF_AW_CHAN_T(aw_chan_t, addr_t, id_t, user_t)
  `AXI_TYPEDEF_W_CHAN_T(mst_w_chan_t, mst_data_t, mst_strb_t, user_t)
  `AXI_TYPEDEF_W_CHAN_T(slv_w_chan_t, slv_data_t, slv_strb_t, user_t)
  `AXI_TYPEDEF_B_CHAN_T(b_chan_t, id_t, user_t)
  `AXI_TYPEDEF_AR_CHAN_T(ar_chan_t, addr_t, id_t, user_t)
  `AXI_TYPEDEF_R_CHAN_T(mst_r_chan_t, mst_data_t, id_t, user_t)
  `AXI_TYPEDEF_R_CHAN_T(slv_r_chan_t, slv_data_t, id_t, user_t)
  `AXI_TYPEDEF_REQ_T(mst_req_t, aw_chan_t, mst_w_chan_t, ar_chan_t)
  `AXI_TYPEDEF_RESP_T(mst_resp_t, b_chan_t, mst_r_chan_t)
  `AXI_TYPEDEF_REQ_T(slv_req_t, aw_chan_t, slv_w_chan_t, ar_chan_t)
  `AXI_TYPEDEF_RESP_T(slv_resp_t, b_chan_t, slv_r_chan_t)

   slv_req_t  axi_req32; 
   slv_resp_t axi_rsp32;
   
   
  // Struct breakout module tool-inserted DFT TAP signals
  pinmux_jtag_breakout u_dft_tap_breakout (
    .req_i    (pinmux_aon_dft_jtag_req),
    .rsp_o    (pinmux_aon_dft_jtag_rsp),
    .tck_o    (),
    .trst_no  (),
    .tms_o    (),
    .tdi_o    (),
    .tdo_i    (1'b0),
    .tdo_oe_i (1'b0)
  );

  simulator_ctrl #(
    .LogName("log.log")
    ) u_simulator_ctrl (
      .clk_i     (clk_main_i),
      .rst_ni    (por_n_i),

      .req_i     (device_req),
      .we_i      (device_we),
      .be_i      (device_be),
      .addr_i    (device_addr),
      .wdata_i   (device_wdata),
      .rvalid_o  (device_rvalid),
      .rdata_o   (device_rdata)

    );
  /* 
  ram_2p #(
      .Depth(1024*1024/4),
      .MemInitFile(SRAMInitFile)
    ) u_ram (
      .clk_i       (clk_main_i),
      .rst_ni      (por_n_i),

      .a_req_i     (device_req[Ram]),
      .a_we_i      (device_we[Ram]),
      .a_be_i      (device_be[Ram]),
      .a_addr_i    (device_addr[Ram]),
      .a_wdata_i   (device_wdata[Ram]),
      .a_rvalid_o  (device_rvalid[Ram]),
      .a_rdata_o   (device_rdata[Ram]),

      .b_req_i     (instr_req),
      .b_we_i      (1'b0),
      .b_be_i      (4'b0),
      .b_addr_i    (instr_addr),
      .b_wdata_i   (32'b0),
      .b_rvalid_o  (instr_rvalid),
      .b_rdata_o   (instr_rdata)
    );*/
   
  axi_dw_converter #(
     .AxiMaxReads        ( AXI_MAX_READS           ),
     .AxiSlvPortDataWidth( AXI_SLV_PORT_DATA_WIDTH ),
     .AxiMstPortDataWidth( AXI_MST_PORT_DATA_WIDTH ),
     .AxiAddrWidth       ( AXI_ADDR_WIDTH          ),
     .AxiIdWidth         ( AXI_ID_WIDTH            ),
     .aw_chan_t          ( aw_chan_t               ),
     .mst_w_chan_t       ( mst_w_chan_t            ),
     .slv_w_chan_t       ( slv_w_chan_t            ),
     .b_chan_t           ( b_chan_t                ),
     .ar_chan_t          ( ar_chan_t               ),
     .mst_r_chan_t       ( mst_r_chan_t            ),
     .slv_r_chan_t       ( slv_r_chan_t            ),
     .axi_mst_req_t      ( mst_req_t               ),
     .axi_mst_resp_t     ( mst_resp_t              ),
     .axi_slv_req_t      ( slv_req_t               ),
     .axi_slv_resp_t     ( slv_resp_t              )
  ) i_axi_dw_converter (
    .clk_i      ( clkmgr_aon_clocks.clk_main_infra    ),
    .rst_ni     ( rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel]   ),
    // slave port
    .slv_req_i  ( axi_req32  ),
    .slv_resp_o ( axi_rsp32  ),
    // master port
    .mst_req_o  ( axi_req  ),
    .mst_resp_i ( axi_rsp  )
  );
   
  tlul2axi #(
      .axi_req_t (slv_req_t),
      .axi_resp_t(slv_resp_t)
  ) u_axi_xbar_mst (
      .rst_ni(rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel]),
      .clk_i(clkmgr_aon_clocks.clk_main_infra),
      .tl_req(core2alsaqr),
      .tl_rsp(alsaqr2core),
      .axi_req(axi_req32),
      .axi_rsp(axi_rsp32)
  );

   assert property (@(posedge axi_req32.w_valid) (core2alsaqr.a_data == axi_req32.w.data));
   assert property (@(posedge axi_req32.r_valid) (alsaqr2core.d_data == axi_rsp32.r.data));

  uart #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[0:0])
  ) u_uart0 (

      // Input
      .cio_rx_i    (cio_uart0_rx_p2d),

      // Output
      .cio_tx_o    (cio_uart0_tx_d2p),
      .cio_tx_en_o (cio_uart0_tx_en_d2p),

      // Interrupt
      .intr_tx_watermark_o  (intr_uart0_tx_watermark),
      .intr_rx_watermark_o  (intr_uart0_rx_watermark),
      .intr_tx_empty_o      (intr_uart0_tx_empty),
      .intr_rx_overflow_o   (intr_uart0_rx_overflow),
      .intr_rx_frame_err_o  (intr_uart0_rx_frame_err),
      .intr_rx_break_err_o  (intr_uart0_rx_break_err),
      .intr_rx_timeout_o    (intr_uart0_rx_timeout),
      .intr_rx_parity_err_o (intr_uart0_rx_parity_err),
      // [0]: fatal_fault
      .alert_tx_o  ( alert_tx[0] ),
      .alert_rx_i  ( alert_rx[0] ),

      // Inter-module signals
      .tl_i(uart0_tl_req),
      .tl_o(uart0_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_peri),
      .rst_ni (rstmgr_aon_resets.rst_sys_io_div4_n[rstmgr_pkg::Domain0Sel])
  );

  uart #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[1:1])
  ) u_uart1 (

      // Input
      .cio_rx_i    (cio_uart1_rx_p2d),

      // Output
      .cio_tx_o    (cio_uart1_tx_d2p),
      .cio_tx_en_o (cio_uart1_tx_en_d2p),

      // Interrupt
      .intr_tx_watermark_o  (intr_uart1_tx_watermark),
      .intr_rx_watermark_o  (intr_uart1_rx_watermark),
      .intr_tx_empty_o      (intr_uart1_tx_empty),
      .intr_rx_overflow_o   (intr_uart1_rx_overflow),
      .intr_rx_frame_err_o  (intr_uart1_rx_frame_err),
      .intr_rx_break_err_o  (intr_uart1_rx_break_err),
      .intr_rx_timeout_o    (intr_uart1_rx_timeout),
      .intr_rx_parity_err_o (intr_uart1_rx_parity_err),
      // [1]: fatal_fault
      .alert_tx_o  ( alert_tx[1:1] ),
      .alert_rx_i  ( alert_rx[1:1] ),

      // Inter-module signals
      .tl_i(uart1_tl_req),
      .tl_o(uart1_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_peri),
      .rst_ni (rstmgr_aon_resets.rst_sys_io_div4_n[rstmgr_pkg::Domain0Sel])
  );

  uart #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[2:2])
  ) u_uart2 (

      // Input
      .cio_rx_i    (cio_uart2_rx_p2d),

      // Output
      .cio_tx_o    (cio_uart2_tx_d2p),
      .cio_tx_en_o (cio_uart2_tx_en_d2p),

      // Interrupt
      .intr_tx_watermark_o  (intr_uart2_tx_watermark),
      .intr_rx_watermark_o  (intr_uart2_rx_watermark),
      .intr_tx_empty_o      (intr_uart2_tx_empty),
      .intr_rx_overflow_o   (intr_uart2_rx_overflow),
      .intr_rx_frame_err_o  (intr_uart2_rx_frame_err),
      .intr_rx_break_err_o  (intr_uart2_rx_break_err),
      .intr_rx_timeout_o    (intr_uart2_rx_timeout),
      .intr_rx_parity_err_o (intr_uart2_rx_parity_err),
      // [2]: fatal_fault
      .alert_tx_o  ( alert_tx[2:2] ),
      .alert_rx_i  ( alert_rx[2:2] ),

      // Inter-module signals
      .tl_i(uart2_tl_req),
      .tl_o(uart2_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_peri),
      .rst_ni (rstmgr_aon_resets.rst_sys_io_div4_n[rstmgr_pkg::Domain0Sel])
  );

  uart #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[3:3])
  ) u_uart3 (

      // Input
      .cio_rx_i    (cio_uart3_rx_p2d),

      // Output
      .cio_tx_o    (cio_uart3_tx_d2p),
      .cio_tx_en_o (cio_uart3_tx_en_d2p),

      // Interrupt
      .intr_tx_watermark_o  (intr_uart3_tx_watermark),
      .intr_rx_watermark_o  (intr_uart3_rx_watermark),
      .intr_tx_empty_o      (intr_uart3_tx_empty),
      .intr_rx_overflow_o   (intr_uart3_rx_overflow),
      .intr_rx_frame_err_o  (intr_uart3_rx_frame_err),
      .intr_rx_break_err_o  (intr_uart3_rx_break_err),
      .intr_rx_timeout_o    (intr_uart3_rx_timeout),
      .intr_rx_parity_err_o (intr_uart3_rx_parity_err),
      // [3]: fatal_fault
      .alert_tx_o  ( alert_tx[3:3] ),
      .alert_rx_i  ( alert_rx[3:3] ),

      // Inter-module signals
      .tl_i(uart3_tl_req),
      .tl_o(uart3_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_peri),
      .rst_ni (rstmgr_aon_resets.rst_sys_io_div4_n[rstmgr_pkg::Domain0Sel])
  );

  gpio #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[4:4])
  ) u_gpio (

      // Input
      .cio_gpio_i    (cio_gpio_gpio_p2d),

      // Output
      .cio_gpio_o    (cio_gpio_gpio_d2p),
      .cio_gpio_en_o (cio_gpio_gpio_en_d2p),

      // Interrupt
      .intr_gpio_o (intr_gpio_gpio),
      // [4]: fatal_fault
      .alert_tx_o  ( alert_tx[4] ),
      .alert_rx_i  ( alert_rx[4] ),

      // Inter-module signals
      .tl_i(gpio_tl_req),
      .tl_o(gpio_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_peri),
      .rst_ni (rstmgr_aon_resets.rst_sys_io_div4_n[rstmgr_pkg::Domain0Sel])
  );

  spi_device #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[5:5])
  ) u_spi_device (

      // Input
      .cio_sck_i    (cio_spi_device_sck_p2d),
      .cio_csb_i    (cio_spi_device_csb_p2d),
      .cio_sd_i     (cio_spi_device_sd_p2d),

      // Output
      .cio_sd_o     (cio_spi_device_sd_d2p),
      .cio_sd_en_o  (cio_spi_device_sd_en_d2p),

      // Interrupt
      .intr_rxf_o         (intr_spi_device_rxf),
      .intr_rxlvl_o       (intr_spi_device_rxlvl),
      .intr_txlvl_o       (intr_spi_device_txlvl),
      .intr_rxerr_o       (intr_spi_device_rxerr),
      .intr_rxoverflow_o  (intr_spi_device_rxoverflow),
      .intr_txunderflow_o (intr_spi_device_txunderflow),
      // [5]: fatal_fault
      .alert_tx_o  ( alert_tx[5] ),
      .alert_rx_i  ( alert_rx[5] ),

      // Inter-module signals
      .ram_cfg_i(ast_ram_2p_cfg),
      .passthrough_o(spi_device_passthrough_req),
      .passthrough_i(spi_device_passthrough_rsp),
      .mbist_en_i('0),
      .tl_i(spi_device_tl_req),
      .tl_o(spi_device_tl_rsp),
      .scanmode_i,
      .scan_rst_ni,

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_peri),
      .scan_clk_i (clkmgr_aon_clocks.clk_io_div2_peri),
      .rst_ni (rstmgr_aon_resets.rst_spi_device_n[rstmgr_pkg::Domain0Sel])
  );

  spi_host #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[6:6])
  ) u_spi_host0 (

      // Input
      .cio_sd_i     (cio_spi_host0_sd_p2d),

      // Output
      .cio_sck_o    (cio_spi_host0_sck_d2p),
      .cio_sck_en_o (cio_spi_host0_sck_en_d2p),
      .cio_csb_o    (cio_spi_host0_csb_d2p),
      .cio_csb_en_o (cio_spi_host0_csb_en_d2p),
      .cio_sd_o     (cio_spi_host0_sd_d2p),
      .cio_sd_en_o  (cio_spi_host0_sd_en_d2p),

      // Interrupt
      .intr_error_o     (intr_spi_host0_error),
      .intr_spi_event_o (intr_spi_host0_spi_event),
      // [6]: fatal_fault
      .alert_tx_o  ( alert_tx[6] ),
      .alert_rx_i  ( alert_rx[6] ),

      // Inter-module signals
      .passthrough_i(spi_device_passthrough_req),
      .passthrough_o(spi_device_passthrough_rsp),
      .tl_i(spi_host0_tl_req),
      .tl_o(spi_host0_tl_rsp),
      .scanmode_i,

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_peri),
      .clk_core_i (clkmgr_aon_clocks.clk_io_peri),
      .rst_ni (rstmgr_aon_resets.rst_spi_host0_n[rstmgr_pkg::Domain0Sel]),
      .rst_core_ni (rstmgr_aon_resets.rst_spi_host0_core_n[rstmgr_pkg::Domain0Sel])
  );
/*
  spi_host #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[7:7])
  ) u_spi_host1 (

      // Input
      .cio_sd_i     (cio_spi_host1_sd_p2d),

      // Output
      .cio_sck_o    (cio_spi_host1_sck_d2p),
      .cio_sck_en_o (cio_spi_host1_sck_en_d2p),
      .cio_csb_o    (cio_spi_host1_csb_d2p),
      .cio_csb_en_o (cio_spi_host1_csb_en_d2p),
      .cio_sd_o     (cio_spi_host1_sd_d2p),
      .cio_sd_en_o  (cio_spi_host1_sd_en_d2p),

      // Interrupt
      .intr_error_o     (intr_spi_host1_error),
      .intr_spi_event_o (intr_spi_host1_spi_event),
      // [7]: fatal_fault
      .alert_tx_o  ( alert_tx[7:7] ),
      .alert_rx_i  ( alert_rx[7:7] ),

      // Inter-module signals
      .passthrough_i(spi_device_pkg::PASSTHROUGH_REQ_DEFAULT),
      .passthrough_o(),
      .tl_i(spi_host1_tl_req),
      .tl_o(spi_host1_tl_rsp),
      .scanmode_i,

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_peri),
      .clk_core_i (clkmgr_aon_clocks.clk_io_div2_peri),
      .rst_ni (rstmgr_aon_resets.rst_spi_host1_n[rstmgr_pkg::Domain0Sel]),
      .rst_core_ni (rstmgr_aon_resets.rst_spi_host1_core_n[rstmgr_pkg::Domain0Sel])
  );*/
/*
  i2c #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[8:8])
  ) u_i2c0 (

      // Input
      .cio_sda_i    (cio_i2c0_sda_p2d),
      .cio_scl_i    (cio_i2c0_scl_p2d),

      // Output
      .cio_sda_o    (cio_i2c0_sda_d2p),
      .cio_sda_en_o (cio_i2c0_sda_en_d2p),
      .cio_scl_o    (cio_i2c0_scl_d2p),
      .cio_scl_en_o (cio_i2c0_scl_en_d2p),

      // Interrupt
      .intr_fmt_watermark_o    (intr_i2c0_fmt_watermark),
      .intr_rx_watermark_o     (intr_i2c0_rx_watermark),
      .intr_fmt_overflow_o     (intr_i2c0_fmt_overflow),
      .intr_rx_overflow_o      (intr_i2c0_rx_overflow),
      .intr_nak_o              (intr_i2c0_nak),
      .intr_scl_interference_o (intr_i2c0_scl_interference),
      .intr_sda_interference_o (intr_i2c0_sda_interference),
      .intr_stretch_timeout_o  (intr_i2c0_stretch_timeout),
      .intr_sda_unstable_o     (intr_i2c0_sda_unstable),
      .intr_trans_complete_o   (intr_i2c0_trans_complete),
      .intr_tx_empty_o         (intr_i2c0_tx_empty),
      .intr_tx_nonempty_o      (intr_i2c0_tx_nonempty),
      .intr_tx_overflow_o      (intr_i2c0_tx_overflow),
      .intr_acq_overflow_o     (intr_i2c0_acq_overflow),
      .intr_ack_stop_o         (intr_i2c0_ack_stop),
      .intr_host_timeout_o     (intr_i2c0_host_timeout),
      // [8]: fatal_fault
      .alert_tx_o  ( alert_tx[8:8] ),
      .alert_rx_i  ( alert_rx[8:8] ),

      // Inter-module signals
      .tl_i(i2c0_tl_req),
      .tl_o(i2c0_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_peri),
      .rst_ni (rstmgr_aon_resets.rst_i2c0_n[rstmgr_pkg::Domain0Sel])
  );

  i2c #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[9:9])
  ) u_i2c1 (

      // Input
      .cio_sda_i    (cio_i2c1_sda_p2d),
      .cio_scl_i    (cio_i2c1_scl_p2d),

      // Output
      .cio_sda_o    (cio_i2c1_sda_d2p),
      .cio_sda_en_o (cio_i2c1_sda_en_d2p),
      .cio_scl_o    (cio_i2c1_scl_d2p),
      .cio_scl_en_o (cio_i2c1_scl_en_d2p),

      // Interrupt
      .intr_fmt_watermark_o    (intr_i2c1_fmt_watermark),
      .intr_rx_watermark_o     (intr_i2c1_rx_watermark),
      .intr_fmt_overflow_o     (intr_i2c1_fmt_overflow),
      .intr_rx_overflow_o      (intr_i2c1_rx_overflow),
      .intr_nak_o              (intr_i2c1_nak),
      .intr_scl_interference_o (intr_i2c1_scl_interference),
      .intr_sda_interference_o (intr_i2c1_sda_interference),
      .intr_stretch_timeout_o  (intr_i2c1_stretch_timeout),
      .intr_sda_unstable_o     (intr_i2c1_sda_unstable),
      .intr_trans_complete_o   (intr_i2c1_trans_complete),
      .intr_tx_empty_o         (intr_i2c1_tx_empty),
      .intr_tx_nonempty_o      (intr_i2c1_tx_nonempty),
      .intr_tx_overflow_o      (intr_i2c1_tx_overflow),
      .intr_acq_overflow_o     (intr_i2c1_acq_overflow),
      .intr_ack_stop_o         (intr_i2c1_ack_stop),
      .intr_host_timeout_o     (intr_i2c1_host_timeout),
      // [9]: fatal_fault
      .alert_tx_o  ( alert_tx[9:9] ),
      .alert_rx_i  ( alert_rx[9:9] ),

      // Inter-module signals
      .tl_i(i2c1_tl_req),
      .tl_o(i2c1_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_peri),
      .rst_ni (rstmgr_aon_resets.rst_i2c1_n[rstmgr_pkg::Domain0Sel])
  );

  i2c #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[10:10])
  ) u_i2c2 (

      // Input
      .cio_sda_i    (cio_i2c2_sda_p2d),
      .cio_scl_i    (cio_i2c2_scl_p2d),

      // Output
      .cio_sda_o    (cio_i2c2_sda_d2p),
      .cio_sda_en_o (cio_i2c2_sda_en_d2p),
      .cio_scl_o    (cio_i2c2_scl_d2p),
      .cio_scl_en_o (cio_i2c2_scl_en_d2p),

      // Interrupt
      .intr_fmt_watermark_o    (intr_i2c2_fmt_watermark),
      .intr_rx_watermark_o     (intr_i2c2_rx_watermark),
      .intr_fmt_overflow_o     (intr_i2c2_fmt_overflow),
      .intr_rx_overflow_o      (intr_i2c2_rx_overflow),
      .intr_nak_o              (intr_i2c2_nak),
      .intr_scl_interference_o (intr_i2c2_scl_interference),
      .intr_sda_interference_o (intr_i2c2_sda_interference),
      .intr_stretch_timeout_o  (intr_i2c2_stretch_timeout),
      .intr_sda_unstable_o     (intr_i2c2_sda_unstable),
      .intr_trans_complete_o   (intr_i2c2_trans_complete),
      .intr_tx_empty_o         (intr_i2c2_tx_empty),
      .intr_tx_nonempty_o      (intr_i2c2_tx_nonempty),
      .intr_tx_overflow_o      (intr_i2c2_tx_overflow),
      .intr_acq_overflow_o     (intr_i2c2_acq_overflow),
      .intr_ack_stop_o         (intr_i2c2_ack_stop),
      .intr_host_timeout_o     (intr_i2c2_host_timeout),
      // [10]: fatal_fault
      .alert_tx_o  ( alert_tx[10:10] ),
      .alert_rx_i  ( alert_rx[10:10] ),

      // Inter-module signals
      .tl_i(i2c2_tl_req),
      .tl_o(i2c2_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_peri),
      .rst_ni (rstmgr_aon_resets.rst_i2c2_n[rstmgr_pkg::Domain0Sel])
  );

  pattgen #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[11:11])
  ) u_pattgen (

      // Output
      .cio_pda0_tx_o    (cio_pattgen_pda0_tx_d2p),
      .cio_pda0_tx_en_o (cio_pattgen_pda0_tx_en_d2p),
      .cio_pcl0_tx_o    (cio_pattgen_pcl0_tx_d2p),
      .cio_pcl0_tx_en_o (cio_pattgen_pcl0_tx_en_d2p),
      .cio_pda1_tx_o    (cio_pattgen_pda1_tx_d2p),
      .cio_pda1_tx_en_o (cio_pattgen_pda1_tx_en_d2p),
      .cio_pcl1_tx_o    (cio_pattgen_pcl1_tx_d2p),
      .cio_pcl1_tx_en_o (cio_pattgen_pcl1_tx_en_d2p),

      // Interrupt
      .intr_done_ch0_o (intr_pattgen_done_ch0),
      .intr_done_ch1_o (intr_pattgen_done_ch1),
      // [11]: fatal_fault
      .alert_tx_o  ( alert_tx[11:11] ),
      .alert_rx_i  ( alert_rx[11:11] ),

      // Inter-module signals
      .tl_i(pattgen_tl_req),
      .tl_o(pattgen_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_peri),
      .rst_ni (rstmgr_aon_resets.rst_sys_io_div4_n[rstmgr_pkg::Domain0Sel])
  );*/

  rv_timer #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[12:12])
  ) u_rv_timer (

      // Interrupt
      .intr_timer_expired_0_0_o (intr_rv_timer_timer_expired_0_0),
      // [12]: fatal_fault
      .alert_tx_o  ( alert_tx[12] ),
      .alert_rx_i  ( alert_rx[12] ),

      // Inter-module signals
      .tl_i(rv_timer_tl_req),
      .tl_o(rv_timer_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_timers),
      .rst_ni (rstmgr_aon_resets.rst_sys_io_div4_n[rstmgr_pkg::Domain0Sel])
  );
/*
  usbdev #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[13:13])
  ) u_usbdev (

      // Input
      .cio_sense_i         (cio_usbdev_sense_p2d),
      .cio_d_i             (cio_usbdev_d_p2d),
      .cio_dp_i            (cio_usbdev_dp_p2d),
      .cio_dn_i            (cio_usbdev_dn_p2d),

      // Output
      .cio_se0_o           (cio_usbdev_se0_d2p),
      .cio_se0_en_o        (cio_usbdev_se0_en_d2p),
      .cio_dp_pullup_o     (cio_usbdev_dp_pullup_d2p),
      .cio_dp_pullup_en_o  (cio_usbdev_dp_pullup_en_d2p),
      .cio_dn_pullup_o     (cio_usbdev_dn_pullup_d2p),
      .cio_dn_pullup_en_o  (cio_usbdev_dn_pullup_en_d2p),
      .cio_tx_mode_se_o    (cio_usbdev_tx_mode_se_d2p),
      .cio_tx_mode_se_en_o (cio_usbdev_tx_mode_se_en_d2p),
      .cio_suspend_o       (cio_usbdev_suspend_d2p),
      .cio_suspend_en_o    (cio_usbdev_suspend_en_d2p),
      .cio_rx_enable_o     (cio_usbdev_rx_enable_d2p),
      .cio_rx_enable_en_o  (cio_usbdev_rx_enable_en_d2p),
      .cio_d_o             (cio_usbdev_d_d2p),
      .cio_d_en_o          (cio_usbdev_d_en_d2p),
      .cio_dp_o            (cio_usbdev_dp_d2p),
      .cio_dp_en_o         (cio_usbdev_dp_en_d2p),
      .cio_dn_o            (cio_usbdev_dn_d2p),
      .cio_dn_en_o         (cio_usbdev_dn_en_d2p),

      // Interrupt
      .intr_pkt_received_o    (intr_usbdev_pkt_received),
      .intr_pkt_sent_o        (intr_usbdev_pkt_sent),
      .intr_disconnected_o    (intr_usbdev_disconnected),
      .intr_host_lost_o       (intr_usbdev_host_lost),
      .intr_link_reset_o      (intr_usbdev_link_reset),
      .intr_link_suspend_o    (intr_usbdev_link_suspend),
      .intr_link_resume_o     (intr_usbdev_link_resume),
      .intr_av_empty_o        (intr_usbdev_av_empty),
      .intr_rx_full_o         (intr_usbdev_rx_full),
      .intr_av_overflow_o     (intr_usbdev_av_overflow),
      .intr_link_in_err_o     (intr_usbdev_link_in_err),
      .intr_rx_crc_err_o      (intr_usbdev_rx_crc_err),
      .intr_rx_pid_err_o      (intr_usbdev_rx_pid_err),
      .intr_rx_bitstuff_err_o (intr_usbdev_rx_bitstuff_err),
      .intr_frame_o           (intr_usbdev_frame),
      .intr_connected_o       (intr_usbdev_connected),
      .intr_link_out_err_o    (intr_usbdev_link_out_err),
      // [13]: fatal_fault
      .alert_tx_o  ( alert_tx[13:13] ),
      .alert_rx_i  ( alert_rx[13:13] ),

      // Inter-module signals
      .usb_ref_val_o(usbdev_usb_ref_val_o),
      .usb_ref_pulse_o(usbdev_usb_ref_pulse_o),
      .usb_out_of_rst_o(usbdev_usb_out_of_rst),
      .usb_aon_wake_en_o(usbdev_usb_aon_wake_en),
      .usb_aon_wake_ack_o(usbdev_usb_aon_wake_ack),
      .usb_suspend_o(usbdev_usb_suspend),
      .usb_state_debug_i(pinmux_aon_usb_state_debug),
      .ram_cfg_i(ast_ram_2p_cfg),
      .tl_i(usbdev_tl_req),
      .tl_o(usbdev_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_peri),
      .clk_aon_i (clkmgr_aon_clocks.clk_aon_peri),
      .clk_usb_48mhz_i (clkmgr_aon_clocks.clk_usb_peri),
      .rst_ni (rstmgr_aon_resets.rst_usb_n[rstmgr_pkg::Domain0Sel]),
      .rst_aon_ni (rstmgr_aon_resets.rst_sys_aon_n[rstmgr_pkg::Domain0Sel]),
      .rst_usb_48mhz_ni (rstmgr_aon_resets.rst_usbif_n[rstmgr_pkg::Domain0Sel])
  );*/

  otp_ctrl #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[16:14]),
    .MemInitFile(OtpCtrlMemInitFile),
    .RndCnstLfsrSeed(RndCnstOtpCtrlLfsrSeed),
    .RndCnstLfsrPerm(RndCnstOtpCtrlLfsrPerm)
  ) u_otp_ctrl (

      // Output
      .cio_test_o    (cio_otp_ctrl_test_d2p),
      .cio_test_en_o (cio_otp_ctrl_test_en_d2p),

      // Interrupt
      .intr_otp_operation_done_o (intr_otp_ctrl_otp_operation_done),
      .intr_otp_error_o          (intr_otp_ctrl_otp_error),
      // [14]: fatal_macro_error
      // [15]: fatal_check_error
      // [16]: fatal_bus_integ_error
      .alert_tx_o  ( alert_tx[16:14] ),
      .alert_rx_i  ( alert_rx[16:14] ),

      // Inter-module signals
      .otp_ext_voltage_h_io(otp_ext_voltage_h_io),
      .otp_ast_pwr_seq_o(otp_ctrl_otp_ast_pwr_seq_o),
      .otp_ast_pwr_seq_h_i(otp_ctrl_otp_ast_pwr_seq_h_i),
      .otp_alert_o(otp_alert_o),
      .edn_o(edn0_edn_req[1]),
      .edn_i(edn0_edn_rsp[1]),
      .pwr_otp_i(pwrmgr_aon_pwr_otp_req),
      .pwr_otp_o(pwrmgr_aon_pwr_otp_rsp),
      .lc_otp_vendor_test_i(lc_ctrl_lc_otp_vendor_test_req),
      .lc_otp_vendor_test_o(lc_ctrl_lc_otp_vendor_test_rsp),
      .lc_otp_program_i(lc_ctrl_lc_otp_program_req),
      .lc_otp_program_o(lc_ctrl_lc_otp_program_rsp),
      .otp_lc_data_o(otp_ctrl_otp_lc_data),
      .lc_escalate_en_i(lc_ctrl_lc_escalate_en),
      .lc_creator_seed_sw_rw_en_i(lc_ctrl_lc_creator_seed_sw_rw_en),
      .lc_seed_hw_rd_en_i(lc_ctrl_lc_seed_hw_rd_en),
      .lc_dft_en_i(lc_ctrl_lc_dft_en),
      .lc_check_byp_en_i(lc_ctrl_lc_check_byp_en),
      .otp_keymgr_key_o(otp_ctrl_otp_keymgr_key),
      .flash_otp_key_i(flash_ctrl_otp_req),
      .flash_otp_key_o(flash_ctrl_otp_rsp),
      .sram_otp_key_i(otp_ctrl_sram_otp_key_req),
      .sram_otp_key_o(otp_ctrl_sram_otp_key_rsp),
      .otbn_otp_key_i(otp_ctrl_otbn_otp_key_req),
      .otbn_otp_key_o(otp_ctrl_otbn_otp_key_rsp),
      .otp_hw_cfg_o(otp_ctrl_otp_hw_cfg),
      .core_tl_i(otp_ctrl_core_tl_req),
      .core_tl_o(otp_ctrl_core_tl_rsp),
      .prim_tl_i(otp_ctrl_prim_tl_req),
      .prim_tl_o(otp_ctrl_prim_tl_rsp),
      .scanmode_i,
      .scan_rst_ni,
      .scan_en_i,

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_secure),
      .clk_edn_i (clkmgr_aon_clocks.clk_main_secure),
      .rst_ni (rstmgr_aon_resets.rst_lc_io_div4_n[rstmgr_pkg::Domain0Sel]),
      .rst_edn_ni (rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel])
  );

  lc_ctrl #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[19:17]),
    .RndCnstLcKeymgrDivInvalid(RndCnstLcCtrlLcKeymgrDivInvalid),
    .RndCnstLcKeymgrDivTestDevRma(RndCnstLcCtrlLcKeymgrDivTestDevRma),
    .RndCnstLcKeymgrDivProduction(RndCnstLcCtrlLcKeymgrDivProduction)
  ) u_lc_ctrl (
      // [17]: fatal_prog_error
      // [18]: fatal_state_error
      // [19]: fatal_bus_integ_error
      .alert_tx_o  ( alert_tx[19:17] ),
      .alert_rx_i  ( alert_rx[19:17] ),

      // Inter-module signals
      .jtag_i(pinmux_aon_lc_jtag_req),
      .jtag_o(pinmux_aon_lc_jtag_rsp),
      .esc_scrap_state0_tx_i(alert_handler_esc_tx[1]),
      .esc_scrap_state0_rx_o(alert_handler_esc_rx[1]),
      .esc_scrap_state1_tx_i(alert_handler_esc_tx[2]),
      .esc_scrap_state1_rx_o(alert_handler_esc_rx[2]),
      .pwr_lc_i(pwrmgr_aon_pwr_lc_req),
      .pwr_lc_o(pwrmgr_aon_pwr_lc_rsp),
      .lc_otp_vendor_test_o(lc_ctrl_lc_otp_vendor_test_req),
      .lc_otp_vendor_test_i(lc_ctrl_lc_otp_vendor_test_rsp),
      .otp_lc_data_i(otp_ctrl_otp_lc_data),
      .lc_otp_program_o(lc_ctrl_lc_otp_program_req),
      .lc_otp_program_i(lc_ctrl_lc_otp_program_rsp),
      .kmac_data_o(kmac_app_req[1]),
      .kmac_data_i(kmac_app_rsp[1]),
      .lc_dft_en_o(lc_ctrl_lc_dft_en),
      .lc_nvm_debug_en_o(lc_ctrl_lc_nvm_debug_en),
      .lc_hw_debug_en_o(lc_ctrl_lc_hw_debug_en),
      .lc_cpu_en_o(lc_ctrl_lc_cpu_en),
      .lc_keymgr_en_o(lc_ctrl_lc_keymgr_en),
      .lc_escalate_en_o(lc_ctrl_lc_escalate_en),
      .lc_clk_byp_req_o(lc_ctrl_lc_clk_byp_req),
      .lc_clk_byp_ack_i(lc_ctrl_lc_clk_byp_ack),
      .lc_flash_rma_req_o(flash_ctrl_rma_req),
      .lc_flash_rma_seed_o(flash_ctrl_rma_seed),
      .lc_flash_rma_ack_i(flash_ctrl_rma_ack),
      .lc_check_byp_en_o(lc_ctrl_lc_check_byp_en),
      .lc_creator_seed_sw_rw_en_o(lc_ctrl_lc_creator_seed_sw_rw_en),
      .lc_owner_seed_sw_rw_en_o(lc_ctrl_lc_owner_seed_sw_rw_en),
      .lc_iso_part_sw_rd_en_o(lc_ctrl_lc_iso_part_sw_rd_en),
      .lc_iso_part_sw_wr_en_o(lc_ctrl_lc_iso_part_sw_wr_en),
      .lc_seed_hw_rd_en_o(lc_ctrl_lc_seed_hw_rd_en),
      .lc_keymgr_div_o(lc_ctrl_lc_keymgr_div),
      .otp_device_id_i(lc_ctrl_otp_device_id),
      .otp_manuf_state_i(lc_ctrl_otp_manuf_state),
      .tl_i(lc_ctrl_tl_req),
      .tl_o(lc_ctrl_tl_rsp),
      .scanmode_i,
      .scan_rst_ni,

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_secure),
      .clk_kmac_i (clkmgr_aon_clocks.clk_main_secure),
      .rst_ni (rstmgr_aon_resets.rst_lc_io_div4_n[rstmgr_pkg::Domain0Sel]),
      .rst_kmac_ni (rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel])
  );

  alert_handler #(
    .RndCnstLfsrSeed(RndCnstAlertHandlerLfsrSeed),
    .RndCnstLfsrPerm(RndCnstAlertHandlerLfsrPerm)
  ) u_alert_handler (

      // Interrupt
      .intr_classa_o (intr_alert_handler_classa),
      .intr_classb_o (intr_alert_handler_classb),
      .intr_classc_o (intr_alert_handler_classc),
      .intr_classd_o (intr_alert_handler_classd),

      // Inter-module signals
      .crashdump_o(alert_handler_crashdump),
      .edn_o(edn0_edn_req[4]),
      .edn_i(edn0_edn_rsp[4]),
      .esc_rx_i(alert_handler_esc_rx),
      .esc_tx_o(alert_handler_esc_tx),
      .tl_i(alert_handler_tl_req),
      .tl_o(alert_handler_tl_rsp),
      // alert signals
      .alert_rx_o  ( alert_rx ),
      .alert_tx_i  ( alert_tx ),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_secure),
      .clk_edn_i (clkmgr_aon_clocks.clk_main_secure),
      .rst_shadowed_ni (rstmgr_aon_resets.rst_lc_io_div4_shadowed_n[rstmgr_pkg::Domain0Sel]),
      .rst_ni (rstmgr_aon_resets.rst_lc_io_div4_n[rstmgr_pkg::Domain0Sel]),
      .rst_edn_ni (rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel])
  );

  pwrmgr #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[20:20])
  ) u_pwrmgr_aon (

      // Interrupt
      .intr_wakeup_o (intr_pwrmgr_aon_wakeup),
      // [20]: fatal_fault
      .alert_tx_o  ( alert_tx[20] ),
      .alert_rx_i  ( alert_rx[20] ),

      // Inter-module signals
      .pwr_ast_o(pwrmgr_ast_req_o),
      .pwr_ast_i(pwrmgr_ast_rsp_i),
      .pwr_rst_o(pwrmgr_aon_pwr_rst_req),
      .pwr_rst_i(pwrmgr_aon_pwr_rst_rsp),
      .pwr_clk_o(pwrmgr_aon_pwr_clk_req),
      .pwr_clk_i(pwrmgr_aon_pwr_clk_rsp),
      .pwr_otp_o(pwrmgr_aon_pwr_otp_req),
      .pwr_otp_i(pwrmgr_aon_pwr_otp_rsp),
      .pwr_lc_o(pwrmgr_aon_pwr_lc_req),
      .pwr_lc_i(pwrmgr_aon_pwr_lc_rsp),
      .pwr_flash_i(pwrmgr_aon_pwr_flash),
      .esc_rst_tx_i(alert_handler_esc_tx[3]),
      .esc_rst_rx_o(alert_handler_esc_rx[3]),
      .pwr_cpu_i(rv_core_ibex_pwrmgr),
      .wakeups_i(pwrmgr_aon_wakeups),
      .rstreqs_i(pwrmgr_aon_rstreqs),
      .strap_o(pwrmgr_aon_strap),

      .low_power_o(pwrmgr_aon_low_power),
      .rom_ctrl_i(rom_ctrl_pwrmgr_data),
      .fetch_en_o(pwrmgr_aon_fetch_en),
      .tl_i(pwrmgr_aon_tl_req),
      .tl_o(pwrmgr_aon_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_powerup),
      .clk_slow_i (clkmgr_aon_clocks.clk_aon_powerup),
      .rst_ni (rstmgr_aon_resets.rst_por_io_div4_n[rstmgr_pkg::DomainAonSel]),
      .rst_slow_ni (rstmgr_aon_resets.rst_por_aon_n[rstmgr_pkg::DomainAonSel])
  );

  rstmgr #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[21:21])
  ) u_rstmgr_aon (
      // [21]: fatal_fault
      .alert_tx_o  ( alert_tx[21] ),
      .alert_rx_i  ( alert_rx[21] ),

      // Inter-module signals
      .por_n_i(por_n_i),
      .pwr_i(pwrmgr_aon_pwr_rst_req),
      .pwr_o(pwrmgr_aon_pwr_rst_rsp),
      .resets_o(rstmgr_aon_resets),
      .rst_cpu_n_i(rv_core_ibex_rst_cpu_n),
      .ndmreset_req_i(rv_dm_ndmreset_req),
      .alert_dump_i(alert_handler_crashdump),
      .cpu_dump_i(rv_core_ibex_crash_dump),
      .resets_ast_o(rsts_ast_o),
      .tl_i(rstmgr_aon_tl_req),
      .tl_o(rstmgr_aon_tl_rsp),
      .scanmode_i,
      .scan_rst_ni,

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_powerup),
      .clk_aon_i (clkmgr_aon_clocks.clk_aon_powerup),
      .clk_main_i (clkmgr_aon_clocks.clk_main_powerup),
      .clk_io_i (clkmgr_aon_clocks.clk_io_powerup),
      .clk_usb_i (clkmgr_aon_clocks.clk_usb_powerup),
      .clk_io_div2_i (clkmgr_aon_clocks.clk_io_div2_powerup),
      .clk_io_div4_i (clkmgr_aon_clocks.clk_io_div4_powerup),
      .rst_ni (rstmgr_aon_resets.rst_por_io_div4_n[rstmgr_pkg::DomainAonSel])
  );

  clkmgr #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[22:22])
  ) u_clkmgr_aon (
      // [22]: fatal_fault
      .alert_tx_o  ( alert_tx[22] ),
      .alert_rx_i  ( alert_rx[22] ),

      // Inter-module signals
      .clocks_o(clkmgr_aon_clocks),
      .lc_dft_en_i(lc_ctrl_lc_dft_en),
      .ast_clk_byp_req_o(ast_clk_byp_req_o),
      .ast_clk_byp_ack_i(ast_clk_byp_ack_i),
      .lc_clk_byp_req_i(lc_ctrl_lc_clk_byp_req),
      .lc_clk_byp_ack_o(lc_ctrl_lc_clk_byp_ack),
      .jitter_en_o(clk_main_jitter_en_o),
      .clk_main_i(clk_main_i),
      .clk_io_i(clk_io_i),
      .clk_usb_i(clk_usb_i),
      .clk_aon_i(clk_aon_i),
      .clocks_ast_o(clks_ast_o),
      .pwr_i(pwrmgr_aon_pwr_clk_req),
      .pwr_o(pwrmgr_aon_pwr_clk_rsp),
      .idle_i(clkmgr_aon_idle),
      .tl_i(clkmgr_aon_tl_req),
      .tl_o(clkmgr_aon_tl_rsp),
      .scanmode_i,

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_powerup),
      .rst_ni (rstmgr_aon_resets.rst_por_io_div4_n[rstmgr_pkg::DomainAonSel]),
      .rst_main_ni (rstmgr_aon_resets.rst_por_n[rstmgr_pkg::DomainAonSel]),
      .rst_io_ni (rstmgr_aon_resets.rst_por_io_n[rstmgr_pkg::DomainAonSel]),
      .rst_usb_ni (rstmgr_aon_resets.rst_por_usb_n[rstmgr_pkg::DomainAonSel]),
      .rst_io_div2_ni (rstmgr_aon_resets.rst_por_io_div2_n[rstmgr_pkg::DomainAonSel]),
      .rst_io_div4_ni (rstmgr_aon_resets.rst_por_io_div4_n[rstmgr_pkg::DomainAonSel])
  );

  sysrst_ctrl #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[23:23])
  ) u_sysrst_ctrl_aon (

      // Input
      .cio_ac_present_i     (cio_sysrst_ctrl_aon_ac_present_p2d),
      .cio_key0_in_i        (cio_sysrst_ctrl_aon_key0_in_p2d),
      .cio_key1_in_i        (cio_sysrst_ctrl_aon_key1_in_p2d),
      .cio_key2_in_i        (cio_sysrst_ctrl_aon_key2_in_p2d),
      .cio_pwrb_in_i        (cio_sysrst_ctrl_aon_pwrb_in_p2d),
      .cio_lid_open_i       (cio_sysrst_ctrl_aon_lid_open_p2d),
      .cio_ec_rst_l_i       (cio_sysrst_ctrl_aon_ec_rst_l_p2d),

      // Output
      .cio_bat_disable_o    (cio_sysrst_ctrl_aon_bat_disable_d2p),
      .cio_bat_disable_en_o (cio_sysrst_ctrl_aon_bat_disable_en_d2p),
      .cio_flash_wp_l_o     (cio_sysrst_ctrl_aon_flash_wp_l_d2p),
      .cio_flash_wp_l_en_o  (cio_sysrst_ctrl_aon_flash_wp_l_en_d2p),
      .cio_key0_out_o       (cio_sysrst_ctrl_aon_key0_out_d2p),
      .cio_key0_out_en_o    (cio_sysrst_ctrl_aon_key0_out_en_d2p),
      .cio_key1_out_o       (cio_sysrst_ctrl_aon_key1_out_d2p),
      .cio_key1_out_en_o    (cio_sysrst_ctrl_aon_key1_out_en_d2p),
      .cio_key2_out_o       (cio_sysrst_ctrl_aon_key2_out_d2p),
      .cio_key2_out_en_o    (cio_sysrst_ctrl_aon_key2_out_en_d2p),
      .cio_pwrb_out_o       (cio_sysrst_ctrl_aon_pwrb_out_d2p),
      .cio_pwrb_out_en_o    (cio_sysrst_ctrl_aon_pwrb_out_en_d2p),
      .cio_z3_wakeup_o      (cio_sysrst_ctrl_aon_z3_wakeup_d2p),
      .cio_z3_wakeup_en_o   (cio_sysrst_ctrl_aon_z3_wakeup_en_d2p),
      .cio_ec_rst_l_o       (cio_sysrst_ctrl_aon_ec_rst_l_d2p),
      .cio_ec_rst_l_en_o    (cio_sysrst_ctrl_aon_ec_rst_l_en_d2p),

      // Interrupt
      .intr_sysrst_ctrl_o (intr_sysrst_ctrl_aon_sysrst_ctrl),
      // [23]: fatal_fault
      .alert_tx_o  ( alert_tx[23] ),
      .alert_rx_i  ( alert_rx[23] ),

      // Inter-module signals
      .aon_sysrst_ctrl_wkup_req_o(pwrmgr_aon_wakeups[0]),
      .aon_sysrst_ctrl_rst_req_o(pwrmgr_aon_rstreqs[0]),
      .tl_i(sysrst_ctrl_aon_tl_req),
      .tl_o(sysrst_ctrl_aon_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_infra),
      .clk_aon_i (clkmgr_aon_clocks.clk_aon_infra),
      .rst_ni (rstmgr_aon_resets.rst_sys_io_div4_n[rstmgr_pkg::DomainAonSel]),
      .rst_aon_ni (rstmgr_aon_resets.rst_sys_aon_n[rstmgr_pkg::DomainAonSel])
  );
/*
  adcctrl #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[24:24])
  ) u_adc_ctrl_aon (

      // Interrupt
      .intr_debug_cable_o (intr_adc_ctrl_aon_debug_cable),
      // [24]: fatal_fault
      .alert_tx_o  ( alert_tx[24:24] ),
      .alert_rx_i  ( alert_rx[24:24] ),

      // Inter-module signals
      .adc_o(adc_req_o),
      .adc_i(adc_rsp_i),
      .debug_cable_wakeup_o(pwrmgr_aon_wakeups[1]),
      .tl_i(adc_ctrl_aon_tl_req),
      .tl_o(adc_ctrl_aon_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_peri),
      .clk_aon_i (clkmgr_aon_clocks.clk_aon_peri),
      .rst_ni (rstmgr_aon_resets.rst_sys_io_div4_n[rstmgr_pkg::DomainAonSel]),
      .rst_aon_ni (rstmgr_aon_resets.rst_sys_aon_n[rstmgr_pkg::DomainAonSel])
  );

  pwm #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[25:25])
  ) u_pwm_aon (

      // Output
      .cio_pwm_o    (cio_pwm_aon_pwm_d2p),
      .cio_pwm_en_o (cio_pwm_aon_pwm_en_d2p),
      // [25]: fatal_fault
      .alert_tx_o  ( alert_tx[25:25] ),
      .alert_rx_i  ( alert_rx[25:25] ),

      // Inter-module signals
      .tl_i(pwm_aon_tl_req),
      .tl_o(pwm_aon_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_powerup),
      .clk_core_i (clkmgr_aon_clocks.clk_aon_powerup),
      .rst_ni (rstmgr_aon_resets.rst_sys_io_div4_n[rstmgr_pkg::DomainAonSel]),
      .rst_core_ni (rstmgr_aon_resets.rst_sys_aon_n[rstmgr_pkg::DomainAonSel])
  );*/
/*
  pinmux #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[26:26]),
    .TargetCfg(PinmuxAonTargetCfg)
  ) u_pinmux_aon (
      // [26]: fatal_fault
      .alert_tx_o  ( alert_tx[26:26] ),
      .alert_rx_i  ( alert_rx[26:26] ),

      // Inter-module signals
      .lc_hw_debug_en_i(lc_ctrl_lc_hw_debug_en),
      .lc_dft_en_i(lc_ctrl_lc_dft_en),
      .lc_jtag_o(pinmux_aon_lc_jtag_req),
      .lc_jtag_i(pinmux_aon_lc_jtag_rsp),
      .rv_jtag_o(pinmux_aon_rv_jtag_req),
      .rv_jtag_i(pinmux_aon_rv_jtag_rsp),
      .dft_jtag_o(pinmux_aon_dft_jtag_req),
      .dft_jtag_i(pinmux_aon_dft_jtag_rsp),
      .dft_strap_test_o(dft_strap_test_o),
      .dft_hold_tap_sel_i(dft_hold_tap_sel_i),
      .sleep_en_i(1'b0),//pwrmgr_aon_low_power),
      .strap_en_i(1'b1),//pwrmgr_aon_strap),
      .aon_wkup_req_o(pwrmgr_aon_wakeups[2]),
      .usb_wkup_req_o(pwrmgr_aon_wakeups[3]),
      .usb_out_of_rst_i(usbdev_usb_out_of_rst),
      .usb_aon_wake_en_i(usbdev_usb_aon_wake_en),
      .usb_aon_wake_ack_i(usbdev_usb_aon_wake_ack),
      .usb_suspend_i(usbdev_usb_suspend),
      .usb_state_debug_o(pinmux_aon_usb_state_debug),
      .tl_i(pinmux_aon_tl_req),
      .tl_o(pinmux_aon_tl_rsp),

      .periph_to_mio_i      (mio_d2p    ),
      .periph_to_mio_oe_i   (mio_en_d2p ),
      .mio_to_periph_o      (mio_p2d    ),

      .mio_attr_o,
      .mio_out_o,
      .mio_oe_o,
      .mio_in_i,

      .periph_to_dio_i      (dio_d2p    ),
      .periph_to_dio_oe_i   (dio_en_d2p ),
      .dio_to_periph_o      (dio_p2d    ),

      .dio_attr_o,
      .dio_out_o,
      .dio_oe_o,
      .dio_in_i,

      .scanmode_i,

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_powerup),
      .clk_aon_i (clkmgr_aon_clocks.clk_aon_powerup),
      .rst_ni (rstmgr_aon_resets.rst_sys_io_div4_n[rstmgr_pkg::DomainAonSel]),
      .rst_aon_ni (rstmgr_aon_resets.rst_sys_aon_n[rstmgr_pkg::DomainAonSel])
  );*/

  aon_timer #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[27:27])
  ) u_aon_timer_aon (

      // Interrupt
      .intr_wkup_timer_expired_o (intr_aon_timer_aon_wkup_timer_expired),
      .intr_wdog_timer_bark_o    (intr_aon_timer_aon_wdog_timer_bark),
      // [27]: fatal_fault
      .alert_tx_o  ( alert_tx[27] ),
      .alert_rx_i  ( alert_rx[27] ),

      // Inter-module signals
      .nmi_wdog_timer_bark_o(aon_timer_aon_nmi_wdog_timer_bark),
      .aon_timer_wkup_req_o(pwrmgr_aon_wakeups[4]),
      .aon_timer_rst_req_o(pwrmgr_aon_rstreqs[1]),
      .lc_escalate_en_i(lc_ctrl_lc_escalate_en),
      .sleep_mode_i(pwrmgr_aon_low_power),
      .tl_i(aon_timer_aon_tl_req),
      .tl_o(aon_timer_aon_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_timers),
      .clk_aon_i (clkmgr_aon_clocks.clk_aon_timers),
      .rst_ni (rstmgr_aon_resets.rst_lc_io_div4_n[rstmgr_pkg::DomainAonSel]),
      .rst_aon_ni (rstmgr_aon_resets.rst_lc_aon_n[rstmgr_pkg::DomainAonSel])
  );
/*
  sensor_ctrl #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[40:28])
  ) u_sensor_ctrl_aon (

      // Output
      .cio_ast_debug_out_o    (cio_sensor_ctrl_aon_ast_debug_out_d2p),
      .cio_ast_debug_out_en_o (cio_sensor_ctrl_aon_ast_debug_out_en_d2p),
      // [28]: recov_as
      // [29]: recov_cg
      // [30]: recov_gd
      // [31]: recov_ts_hi
      // [32]: recov_ts_lo
      // [33]: recov_fla
      // [34]: recov_otp
      // [35]: recov_ot0
      // [36]: recov_ot1
      // [37]: recov_ot2
      // [38]: recov_ot3
      // [39]: recov_ot4
      // [40]: recov_ot5
      .alert_tx_o  ( alert_tx[40:28] ),
      .alert_rx_i  ( alert_rx[40:28] ),

      // Inter-module signals
      .ast_alert_i(sensor_ctrl_ast_alert_req_i),
      .ast_alert_o(sensor_ctrl_ast_alert_rsp_o),
      .ast_status_i(sensor_ctrl_ast_status_i),
      .ast_init_done_i(ast_init_done_i),
      .ast2pinmux_i(ast2pinmux_i),
      .tl_i(sensor_ctrl_aon_tl_req),
      .tl_o(sensor_ctrl_aon_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_secure),
      .rst_ni (rstmgr_aon_resets.rst_lc_io_div4_n[rstmgr_pkg::DomainAonSel])
  );*/

  sram_ctrl #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[41:41]),
    .RndCnstSramKey(RndCnstSramCtrlRetAonSramKey),
    .RndCnstSramNonce(RndCnstSramCtrlRetAonSramNonce),
    .RndCnstLfsrSeed(RndCnstSramCtrlRetAonLfsrSeed),
    .RndCnstLfsrPerm(RndCnstSramCtrlRetAonLfsrPerm),
    .MemSizeRam(4096),
    .InstrExec(SramCtrlRetAonInstrExec)
  ) u_sram_ctrl_ret_aon (
      // [41]: fatal_error
      .alert_tx_o  ( alert_tx[41] ),
      .alert_rx_i  ( alert_rx[41] ),

      // Inter-module signals
      .sram_otp_key_o(otp_ctrl_sram_otp_key_req[1]),
      .sram_otp_key_i(otp_ctrl_sram_otp_key_rsp[1]),
      .cfg_i(ast_ram_1p_cfg),
      .lc_escalate_en_i(lc_ctrl_lc_escalate_en),
      .lc_hw_debug_en_i(lc_ctrl_lc_hw_debug_en),
      .otp_en_sram_ifetch_i('0),
      .regs_tl_i(sram_ctrl_ret_aon_regs_tl_req),
      .regs_tl_o(sram_ctrl_ret_aon_regs_tl_rsp),
      .ram_tl_i(sram_ctrl_ret_aon_ram_tl_req),
      .ram_tl_o(sram_ctrl_ret_aon_ram_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_io_div4_infra),
      .clk_otp_i (clkmgr_aon_clocks.clk_io_div4_infra),
      .rst_ni (rstmgr_aon_resets.rst_sys_io_div4_n[rstmgr_pkg::DomainAonSel]),
      .rst_otp_ni (rstmgr_aon_resets.rst_lc_io_div4_n[rstmgr_pkg::DomainAonSel])
  );

  flash_ctrl #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[45:42]),
    .RndCnstAddrKey(RndCnstFlashCtrlAddrKey),
    .RndCnstDataKey(RndCnstFlashCtrlDataKey),
    .RndCnstLfsrSeed(RndCnstFlashCtrlLfsrSeed),
    .RndCnstLfsrPerm(RndCnstFlashCtrlLfsrPerm)
  ) u_flash_ctrl (

      // Input
      .cio_tck_i    (cio_flash_ctrl_tck_p2d),
      .cio_tms_i    (cio_flash_ctrl_tms_p2d),
      .cio_tdi_i    (cio_flash_ctrl_tdi_p2d),

      // Output
      .cio_tdo_o    (cio_flash_ctrl_tdo_d2p),
      .cio_tdo_en_o (cio_flash_ctrl_tdo_en_d2p),

      // Interrupt
      .intr_prog_empty_o (intr_flash_ctrl_prog_empty),
      .intr_prog_lvl_o   (intr_flash_ctrl_prog_lvl),
      .intr_rd_full_o    (intr_flash_ctrl_rd_full),
      .intr_rd_lvl_o     (intr_flash_ctrl_rd_lvl),
      .intr_op_done_o    (intr_flash_ctrl_op_done),
      .intr_err_o        (intr_flash_ctrl_err),
      // [42]: recov_err
      // [43]: recov_mp_err
      // [44]: recov_ecc_err
      // [45]: fatal_intg_err
      .alert_tx_o  ( alert_tx[45:42] ),
      .alert_rx_i  ( alert_rx[45:42] ),

      // Inter-module signals
      .otp_o(flash_ctrl_otp_req),
      .otp_i(flash_ctrl_otp_rsp),
      .lc_nvm_debug_en_i(lc_ctrl_lc_nvm_debug_en),
      .flash_bist_enable_i(flash_bist_enable_i),
      .flash_power_down_h_i(flash_power_down_h_i),
      .flash_power_ready_h_i(flash_power_ready_h_i),
      .flash_test_mode_a_io(flash_test_mode_a_io),
      .flash_test_voltage_h_io(flash_test_voltage_h_io),
      .flash_alert_o(flash_alert_o),
      .lc_creator_seed_sw_rw_en_i(lc_ctrl_lc_creator_seed_sw_rw_en),
      .lc_owner_seed_sw_rw_en_i(lc_ctrl_lc_owner_seed_sw_rw_en),
      .lc_iso_part_sw_rd_en_i(lc_ctrl_lc_iso_part_sw_rd_en),
      .lc_iso_part_sw_wr_en_i(lc_ctrl_lc_iso_part_sw_wr_en),
      .lc_seed_hw_rd_en_i(lc_ctrl_lc_seed_hw_rd_en),
      .lc_escalate_en_i(lc_ctrl_lc_escalate_en),
      .rma_req_i(flash_ctrl_rma_req),
      .rma_ack_o(flash_ctrl_rma_ack),
      .rma_seed_i(flash_ctrl_rma_seed),
      .pwrmgr_o(pwrmgr_aon_pwr_flash),
      .keymgr_o(flash_ctrl_keymgr),
      .core_tl_i(flash_ctrl_core_tl_req),
      .core_tl_o(flash_ctrl_core_tl_rsp),
      .prim_tl_i(flash_ctrl_prim_tl_req),
      .prim_tl_o(flash_ctrl_prim_tl_rsp),
      .mem_tl_i(flash_ctrl_mem_tl_req),
      .mem_tl_o(flash_ctrl_mem_tl_rsp),
      .scanmode_i,
      .scan_rst_ni,
      .scan_en_i,

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_main_infra),
      .clk_otp_i (clkmgr_aon_clocks.clk_io_div4_infra),
      .rst_ni (rstmgr_aon_resets.rst_lc_n[rstmgr_pkg::Domain0Sel]),
      .rst_otp_ni (rstmgr_aon_resets.rst_lc_io_div4_n[rstmgr_pkg::Domain0Sel])
  );

  rv_dm #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[46:46]),
    .IdcodeValue(RvDmIdcodeValue)
  ) u_rv_dm (
      // [46]: fatal_fault
      .alert_tx_o  ( alert_tx[46] ),
      .alert_rx_i  ( alert_rx[46] ),

      // Inter-module signals
      .jtag_i,//pinmux_aon_rv_jtag_req),
      .jtag_o,//pinmux_aon_rv_jtag_rsp),
      .lc_hw_debug_en_i(lc_ctrl_pkg::On),//lc_ctrl_lc_hw_debug_en),
      .unavailable_i(1'b0),
      .ndmreset_req_o(rv_dm_ndmreset_req),
      .dmactive_o(),
      .debug_req_o(rv_dm_debug_req),
      .sba_tl_h_o(main_tl_rv_dm__sba_req),
      .sba_tl_h_i(main_tl_rv_dm__sba_rsp),
      .regs_tl_d_i(rv_dm_regs_tl_d_req),
      .regs_tl_d_o(rv_dm_regs_tl_d_rsp),
      .rom_tl_d_i(rv_dm_rom_tl_d_req),
      .rom_tl_d_o(rv_dm_rom_tl_d_rsp),
      .scanmode_i,
      .scan_rst_ni,

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_main_infra),
      .rst_ni (rstmgr_aon_resets.rst_lc_n[rstmgr_pkg::Domain0Sel])
  );

  rv_ibex_plic #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[47:47])
  ) u_rv_plic (
      // [47]: fatal_fault
      .alert_tx_o  ( alert_tx[47] ),
      .alert_rx_i  ( alert_rx[47] ),

      // Inter-module signals
      .irq_o(rv_plic_irq),
      .irq_id_o(),
      .msip_o(rv_plic_msip),
      .tl_i(rv_plic_tl_req),
      .tl_o(rv_plic_tl_rsp),
      .intr_src_i (intr_vector),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_main_secure),
      .rst_ni (rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel])
  );

  aes #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[49:48]),
    .AES192Enable(1'b1),
    .Masking(AesMasking),
    .SBoxImpl(AesSBoxImpl),
    .SecStartTriggerDelay(SecAesStartTriggerDelay),
    .SecAllowForcingMasks(SecAesAllowForcingMasks),
    .SecSkipPRNGReseeding(SecAesSkipPRNGReseeding),
    .RndCnstClearingLfsrSeed(RndCnstAesClearingLfsrSeed),
    .RndCnstClearingLfsrPerm(RndCnstAesClearingLfsrPerm),
    .RndCnstClearingSharePerm(RndCnstAesClearingSharePerm),
    .RndCnstMaskingLfsrSeed(RndCnstAesMaskingLfsrSeed),
    .RndCnstMskgChunkLfsrPerm(RndCnstAesMskgChunkLfsrPerm)
  ) u_aes (
      // [48]: recov_ctrl_update_err
      // [49]: fatal_fault
      .alert_tx_o  ( alert_tx[49:48] ),
      .alert_rx_i  ( alert_rx[49:48] ),

      // Inter-module signals
      .idle_o(clkmgr_aon_idle[0]),
      .lc_escalate_en_i(lc_ctrl_lc_escalate_en),
      .edn_o(edn0_edn_req[5]),
      .edn_i(edn0_edn_rsp[5]),
      .tl_i(aes_tl_req),
      .tl_o(aes_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_main_aes),
      .clk_edn_i (clkmgr_aon_clocks.clk_main_aes),
      .rst_shadowed_ni (rstmgr_aon_resets.rst_sys_shadowed_n[rstmgr_pkg::Domain0Sel]),
      .rst_ni (rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel]),
      .rst_edn_ni (rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel])
  );

  hmac #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[50:50])
  ) u_hmac (

      // Interrupt
      .intr_hmac_done_o  (intr_hmac_hmac_done),
      .intr_fifo_empty_o (intr_hmac_fifo_empty),
      .intr_hmac_err_o   (intr_hmac_hmac_err),
      // [50]: fatal_fault
      .alert_tx_o  ( alert_tx[50] ),
      .alert_rx_i  ( alert_rx[50] ),

      // Inter-module signals
      .idle_o(clkmgr_aon_idle[1]),
      .tl_i(hmac_tl_req),
      .tl_o(hmac_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_main_hmac),
      .rst_ni (rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel])
  );

  kmac #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[51:51]),
    .EnMasking(KmacEnMasking),
    .ReuseShare(KmacReuseShare),
    .RndCnstLfsrPerm(RndCnstKmacLfsrPerm)
  ) u_kmac (

      // Interrupt
      .intr_kmac_done_o  (intr_kmac_kmac_done),
      .intr_fifo_empty_o (intr_kmac_fifo_empty),
      .intr_kmac_err_o   (intr_kmac_kmac_err),
      // [51]: fatal_fault
      .alert_tx_o  ( alert_tx[51] ),
      .alert_rx_i  ( alert_rx[51] ),

      // Inter-module signals
      .keymgr_key_i(keymgr_kmac_key),
      .app_i(kmac_app_req),
      .app_o(kmac_app_rsp),
      .entropy_o(edn0_edn_req[3]),
      .entropy_i(edn0_edn_rsp[3]),
      .idle_o(clkmgr_aon_idle[2]),
      .en_masking_o(kmac_en_masking),
      .tl_i(kmac_tl_req),
      .tl_o(kmac_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_main_kmac),
      .clk_edn_i (clkmgr_aon_clocks.clk_main_kmac),
      .rst_ni (rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel]),
      .rst_edn_ni (rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel])
  );

  keymgr #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[53:52]),
    .KmacEnMasking(KeymgrKmacEnMasking),
    .RndCnstLfsrSeed(RndCnstKeymgrLfsrSeed),
    .RndCnstLfsrPerm(RndCnstKeymgrLfsrPerm),
    .RndCnstRandPerm(RndCnstKeymgrRandPerm),
    .RndCnstRevisionSeed(RndCnstKeymgrRevisionSeed),
    .RndCnstCreatorIdentitySeed(RndCnstKeymgrCreatorIdentitySeed),
    .RndCnstOwnerIntIdentitySeed(RndCnstKeymgrOwnerIntIdentitySeed),
    .RndCnstOwnerIdentitySeed(RndCnstKeymgrOwnerIdentitySeed),
    .RndCnstSoftOutputSeed(RndCnstKeymgrSoftOutputSeed),
    .RndCnstHardOutputSeed(RndCnstKeymgrHardOutputSeed),
    .RndCnstAesSeed(RndCnstKeymgrAesSeed),
    .RndCnstKmacSeed(RndCnstKeymgrKmacSeed),
    .RndCnstOtbnSeed(RndCnstKeymgrOtbnSeed),
    .RndCnstNoneSeed(RndCnstKeymgrNoneSeed)
  ) u_keymgr (

      // Interrupt
      .intr_op_done_o (intr_keymgr_op_done),
      // [52]: fatal_fault_err
      // [53]: recov_operation_err
      .alert_tx_o  ( alert_tx[53:52] ),
      .alert_rx_i  ( alert_rx[53:52] ),

      // Inter-module signals
      .edn_o(edn0_edn_req[0]),
      .edn_i(edn0_edn_rsp[0]),
      .aes_key_o(),
      .kmac_key_o(keymgr_kmac_key),
      .otbn_key_o(),
      .kmac_data_o(kmac_app_req[0]),
      .kmac_data_i(kmac_app_rsp[0]),
      .otp_key_i(otp_ctrl_otp_keymgr_key),
      .otp_device_id_i(keymgr_otp_device_id),
      .flash_i(flash_ctrl_keymgr),
      .lc_keymgr_en_i(lc_ctrl_lc_keymgr_en),
      .lc_keymgr_div_i(lc_ctrl_lc_keymgr_div),
      .rom_digest_i(rom_ctrl_keymgr_data),
      .kmac_en_masking_i(kmac_en_masking),
      .tl_i(keymgr_tl_req),
      .tl_o(keymgr_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_main_secure),
      .clk_edn_i (clkmgr_aon_clocks.clk_main_secure),
      .rst_shadowed_ni (rstmgr_aon_resets.rst_sys_shadowed_n[rstmgr_pkg::Domain0Sel]),
      .rst_ni (rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel]),
      .rst_edn_ni (rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel])
  );

  csrng #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[55:54]),
    .RndCnstCsKeymgrDivNonProduction(RndCnstCsrngCsKeymgrDivNonProduction),
    .RndCnstCsKeymgrDivProduction(RndCnstCsrngCsKeymgrDivProduction),
    .SBoxImpl(CsrngSBoxImpl)
  ) u_csrng (

      // Interrupt
      .intr_cs_cmd_req_done_o (intr_csrng_cs_cmd_req_done),
      .intr_cs_entropy_req_o  (intr_csrng_cs_entropy_req),
      .intr_cs_hw_inst_exc_o  (intr_csrng_cs_hw_inst_exc),
      .intr_cs_fatal_err_o    (intr_csrng_cs_fatal_err),
      // [54]: recov_alert
      // [55]: fatal_alert
      .alert_tx_o  ( alert_tx[55:54] ),
      .alert_rx_i  ( alert_rx[55:54] ),

      // Inter-module signals
      .csrng_cmd_i(csrng_csrng_cmd_req),
      .csrng_cmd_o(csrng_csrng_cmd_rsp),
      .entropy_src_hw_if_o(csrng_entropy_src_hw_if_req),
      .entropy_src_hw_if_i(csrng_entropy_src_hw_if_rsp),
      .cs_aes_halt_i(csrng_cs_aes_halt_req),
      .cs_aes_halt_o(csrng_cs_aes_halt_rsp),
      .otp_en_csrng_sw_app_read_i(csrng_otp_en_csrng_sw_app_read),
      .lc_hw_debug_en_i(lc_ctrl_lc_hw_debug_en),
      .tl_i(csrng_tl_req),
      .tl_o(csrng_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_main_secure),
      .rst_ni (rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel])
  );

  entropy_src #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[57:56]),
    .Stub(EntropySrcStub)
  ) u_entropy_src (

      // Interrupt
      .intr_es_entropy_valid_o      (intr_entropy_src_es_entropy_valid),
      .intr_es_health_test_failed_o (intr_entropy_src_es_health_test_failed),
      .intr_es_observe_fifo_ready_o (intr_entropy_src_es_observe_fifo_ready),
      .intr_es_fatal_err_o          (intr_entropy_src_es_fatal_err),
      // [56]: recov_alert
      // [57]: fatal_alert
      .alert_tx_o  ( alert_tx[57:56] ),
      .alert_rx_i  ( alert_rx[57:56] ),

      // Inter-module signals
      .entropy_src_hw_if_i(csrng_entropy_src_hw_if_req),
      .entropy_src_hw_if_o(csrng_entropy_src_hw_if_rsp),
      .cs_aes_halt_o(csrng_cs_aes_halt_req),
      .cs_aes_halt_i(csrng_cs_aes_halt_rsp),
      .entropy_src_rng_o(es_rng_req_o),
      .entropy_src_rng_i(es_rng_rsp_i),
      .entropy_src_xht_o(),
      .entropy_src_xht_i(entropy_src_pkg::ENTROPY_SRC_XHT_RSP_DEFAULT),
      .otp_en_entropy_src_fw_read_i(entropy_src_otp_en_entropy_src_fw_read),
      .otp_en_entropy_src_fw_over_i(entropy_src_otp_en_entropy_src_fw_over),
      .rng_fips_o(es_rng_fips_o),
      .tl_i(entropy_src_tl_req),
      .tl_o(entropy_src_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_main_secure),
      .rst_ni (rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel])
  );

  edn #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[59:58])
  ) u_edn0 (

      // Interrupt
      .intr_edn_cmd_req_done_o (intr_edn0_edn_cmd_req_done),
      .intr_edn_fatal_err_o    (intr_edn0_edn_fatal_err),
      // [58]: recov_alert
      // [59]: fatal_alert
      .alert_tx_o  ( alert_tx[59:58] ),
      .alert_rx_i  ( alert_rx[59:58] ),

      // Inter-module signals
      .csrng_cmd_o(csrng_csrng_cmd_req[0]),
      .csrng_cmd_i(csrng_csrng_cmd_rsp[0]),
      .edn_i(edn0_edn_req),
      .edn_o(edn0_edn_rsp),
      .tl_i(edn0_tl_req),
      .tl_o(edn0_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_main_secure),
      .rst_ni (rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel])
  );

  edn #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[61:60])
  ) u_edn1 (

      // Interrupt
      .intr_edn_cmd_req_done_o (intr_edn1_edn_cmd_req_done),
      .intr_edn_fatal_err_o    (intr_edn1_edn_fatal_err),
      // [60]: recov_alert
      // [61]: fatal_alert
      .alert_tx_o  ( alert_tx[61:60] ),
      .alert_rx_i  ( alert_rx[61:60] ),

      // Inter-module signals
      .csrng_cmd_o(csrng_csrng_cmd_req[1]),
      .csrng_cmd_i(csrng_csrng_cmd_rsp[1]),
      .edn_i(edn1_edn_req),
      .edn_o(edn1_edn_rsp),
      .tl_i(edn1_tl_req),
      .tl_o(edn1_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_main_secure),
      .rst_ni (rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel])
  );

  sram_ctrl #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[62:62]),
    .RndCnstSramKey(RndCnstSramCtrlMainSramKey),
    .RndCnstSramNonce(RndCnstSramCtrlMainSramNonce),
    .RndCnstLfsrSeed(RndCnstSramCtrlMainLfsrSeed),
    .RndCnstLfsrPerm(RndCnstSramCtrlMainLfsrPerm),
    .MemSizeRam(131072),
    .InstrExec(SramCtrlMainInstrExec)
  ) u_sram_ctrl_main (
      // [62]: fatal_error
      .alert_tx_o  ( alert_tx[62] ),
      .alert_rx_i  ( alert_rx[62] ),

      // Inter-module signals
      .sram_otp_key_o(otp_ctrl_sram_otp_key_req[0]),
      .sram_otp_key_i(otp_ctrl_sram_otp_key_rsp[0]),
      .cfg_i(ast_ram_1p_cfg),
      .lc_escalate_en_i(lc_ctrl_lc_escalate_en),
      .lc_hw_debug_en_i(lc_ctrl_lc_hw_debug_en),
      .otp_en_sram_ifetch_i(sram_ctrl_main_otp_en_sram_ifetch),//prim_mubi_pkg::MuBi8True),//
      .regs_tl_i(sram_ctrl_main_regs_tl_req),
      .regs_tl_o(sram_ctrl_main_regs_tl_rsp),
      .ram_tl_i(sram_ctrl_main_ram_tl_req),
      .ram_tl_o(sram_ctrl_main_ram_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_main_infra),
      .clk_otp_i (clkmgr_aon_clocks.clk_io_div4_infra),
      .rst_ni (rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel]),
      .rst_otp_ni (rstmgr_aon_resets.rst_lc_io_div4_n[rstmgr_pkg::Domain0Sel])
  );

  otbn #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[64:63]),
    .Stub(OtbnStub),
    .RegFile(OtbnRegFile),
    .RndCnstUrndLfsrSeed(RndCnstOtbnUrndLfsrSeed),
    .RndCnstUrndChunkLfsrPerm(RndCnstOtbnUrndChunkLfsrPerm),
    .RndCnstOtbnKey(RndCnstOtbnOtbnKey),
    .RndCnstOtbnNonce(RndCnstOtbnOtbnNonce)
  ) u_otbn (

      // Interrupt
      .intr_done_o (intr_otbn_done),
      // [63]: fatal
      // [64]: recov
      .alert_tx_o  ( alert_tx[64:63] ),
      .alert_rx_i  ( alert_rx[64:63] ),

      // Inter-module signals
      .otbn_otp_key_o(otp_ctrl_otbn_otp_key_req),
      .otbn_otp_key_i(otp_ctrl_otbn_otp_key_rsp),
      .edn_rnd_o(edn1_edn_req[0]),
      .edn_rnd_i(edn1_edn_rsp[0]),
      .edn_urnd_o(edn0_edn_req[6]),
      .edn_urnd_i(edn0_edn_rsp[6]),
      .idle_o(clkmgr_aon_idle[4]),
      .idle_otp_o(clkmgr_aon_idle[3]),
      .ram_cfg_i(ast_ram_1p_cfg),
      .lc_escalate_en_i(lc_ctrl_lc_escalate_en),
      .tl_i(otbn_tl_req),
      .tl_o(otbn_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_main_otbn),
      .clk_edn_i (clkmgr_aon_clocks.clk_main_otbn),
      .clk_otp_i (clkmgr_aon_clocks.clk_io_div4_otbn),
      .rst_ni (rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel]),
      .rst_edn_ni (rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel]),
      .rst_otp_ni (rstmgr_aon_resets.rst_lc_io_div4_n[rstmgr_pkg::Domain0Sel])
  );

  rom_ctrl #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[65:65]),
    .BootRomInitFile(RomCtrlBootRomInitFile),
    .RndCnstScrNonce(RndCnstRomCtrlScrNonce),
    .RndCnstScrKey(RndCnstRomCtrlScrKey),
    .SecDisableScrambling(SecRomCtrlDisableScrambling)
  ) u_rom_ctrl (
      // [65]: fatal
      .alert_tx_o  ( alert_tx[65] ),
      .alert_rx_i  ( alert_rx[65] ),

      // Inter-module signals
      .rom_cfg_i(ast_rom_cfg),
      .pwrmgr_data_o(rom_ctrl_pwrmgr_data),
      .keymgr_data_o(rom_ctrl_keymgr_data),
      .kmac_data_o(kmac_app_req[2]),
      .kmac_data_i(kmac_app_rsp[2]),
      .regs_tl_i(rom_ctrl_regs_tl_req),
      .regs_tl_o(rom_ctrl_regs_tl_rsp),
      .rom_tl_i(rom_ctrl_rom_tl_req),
      .rom_tl_o(rom_ctrl_rom_tl_rsp),

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_main_infra),
      .rst_ni (rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel])
  );

  rv_core_ibex #(
    .AlertAsyncOn(alert_handler_reg_pkg::AsyncOn[69:66]),
    .RndCnstLfsrSeed(RndCnstRvCoreIbexLfsrSeed),
    .RndCnstLfsrPerm(RndCnstRvCoreIbexLfsrPerm),
    .PMPEnable(RvCoreIbexPMPEnable),
    .PMPGranularity(RvCoreIbexPMPGranularity),
    .PMPNumRegions(RvCoreIbexPMPNumRegions),
    .MHPMCounterNum(RvCoreIbexMHPMCounterNum),
    .MHPMCounterWidth(RvCoreIbexMHPMCounterWidth),
    .RV32E(RvCoreIbexRV32E),
    .RV32M(RvCoreIbexRV32M),
    .RV32B(RvCoreIbexRV32B),
    .RegFile(RvCoreIbexRegFile),
    .BranchTargetALU(RvCoreIbexBranchTargetALU),
    .WritebackStage(RvCoreIbexWritebackStage),
    .ICache(RvCoreIbexICache),
    .ICacheECC(RvCoreIbexICacheECC),
    .BranchPredictor(RvCoreIbexBranchPredictor),
    .DbgTriggerEn(RvCoreIbexDbgTriggerEn),
    .SecureIbex(RvCoreIbexSecureIbex),
    .DmHaltAddr(RvCoreIbexDmHaltAddr),
    .DmExceptionAddr(RvCoreIbexDmExceptionAddr),
    .PipeLine(RvCoreIbexPipeLine)
  ) u_rv_core_ibex (
      // [66]: fatal_sw_err
      // [67]: recov_sw_err
      // [68]: fatal_hw_err
      // [69]: recov_hw_err
      .alert_tx_o  ( alert_tx[69:66] ),
      .alert_rx_i  ( alert_rx[69:66] ),

      // Inter-module signals
      .rst_cpu_n_o(rv_core_ibex_rst_cpu_n),
      .ram_cfg_i(ast_ram_1p_cfg),
      .hart_id_i(rv_core_ibex_hart_id),
      .boot_addr_i(rv_core_ibex_boot_addr),
      .irq_software_i(rv_plic_msip),
      .irq_timer_i(rv_core_ibex_irq_timer),
      .irq_external_i(rv_plic_irq),
      .esc_tx_i(alert_handler_esc_tx[0]),
      .esc_rx_o(alert_handler_esc_rx[0]),
      .debug_req_i(rv_dm_debug_req),
      .crash_dump_o(rv_core_ibex_crash_dump),
      .lc_cpu_en_i(lc_ctrl_lc_cpu_en),
      .pwrmgr_cpu_en_i(pwrmgr_aon_fetch_en),
      .pwrmgr_o(rv_core_ibex_pwrmgr),
      .nmi_wdog_i(aon_timer_aon_nmi_wdog_timer_bark),
      .corei_tl_h_o(main_tl_rv_core_ibex__corei_req),//core2instr),//
      .corei_tl_h_i(main_tl_rv_core_ibex__corei_rsp),//instr2core),//
      .cored_tl_h_o(main_tl_rv_core_ibex__cored_req),
      .cored_tl_h_i(main_tl_rv_core_ibex__cored_rsp),
      .cfg_tl_d_i(rv_core_ibex_cfg_tl_d_req),
      .cfg_tl_d_o(rv_core_ibex_cfg_tl_d_rsp),
      .scanmode_i,
      .scan_rst_ni,

      // Clock and reset connections
      .clk_i (clkmgr_aon_clocks.clk_main_infra),//clk_main_i),//
      .clk_esc_i (clkmgr_aon_clocks.clk_io_div4_infra),//(clk_main_i),//
      .rst_ni (rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel]),//(por_n_i),//
      .rst_esc_ni (rstmgr_aon_resets.rst_lc_io_div4_n[rstmgr_pkg::Domain0Sel])//(por_n_i)//
  );

  // interrupt assignments
  assign intr_vector = {
      intr_otbn_done, // IDs [179 +: 1]
      intr_edn1_edn_fatal_err, // IDs [178 +: 1]
      intr_edn1_edn_cmd_req_done, // IDs [177 +: 1]
      intr_edn0_edn_fatal_err, // IDs [176 +: 1]
      intr_edn0_edn_cmd_req_done, // IDs [175 +: 1]
      intr_entropy_src_es_fatal_err, // IDs [174 +: 1]
      intr_entropy_src_es_observe_fifo_ready, // IDs [173 +: 1]
      intr_entropy_src_es_health_test_failed, // IDs [172 +: 1]
      intr_entropy_src_es_entropy_valid, // IDs [171 +: 1]
      intr_csrng_cs_fatal_err, // IDs [170 +: 1]
      intr_csrng_cs_hw_inst_exc, // IDs [169 +: 1]
      intr_csrng_cs_entropy_req, // IDs [168 +: 1]
      intr_csrng_cs_cmd_req_done, // IDs [167 +: 1]
      intr_keymgr_op_done, // IDs [166 +: 1]
      intr_kmac_kmac_err, // IDs [165 +: 1]
      intr_kmac_fifo_empty, // IDs [164 +: 1]
      intr_kmac_kmac_done, // IDs [163 +: 1]
      intr_hmac_hmac_err, // IDs [162 +: 1]
      intr_hmac_fifo_empty, // IDs [161 +: 1]
      intr_hmac_hmac_done, // IDs [160 +: 1]
      intr_flash_ctrl_err, // IDs [159 +: 1]
      intr_flash_ctrl_op_done, // IDs [158 +: 1]
      intr_flash_ctrl_rd_lvl, // IDs [157 +: 1]
      intr_flash_ctrl_rd_full, // IDs [156 +: 1]
      intr_flash_ctrl_prog_lvl, // IDs [155 +: 1]
      intr_flash_ctrl_prog_empty, // IDs [154 +: 1]
      intr_aon_timer_aon_wdog_timer_bark, // IDs [153 +: 1]
      intr_aon_timer_aon_wkup_timer_expired, // IDs [152 +: 1]
      1'b0,//intr_adc_ctrl_aon_debug_cable, // IDs [151 +: 1]
      intr_sysrst_ctrl_aon_sysrst_ctrl, // IDs [150 +: 1]
      intr_pwrmgr_aon_wakeup, // IDs [149 +: 1]
      intr_alert_handler_classd, // IDs [148 +: 1]
      intr_alert_handler_classc, // IDs [147 +: 1]
      intr_alert_handler_classb, // IDs [146 +: 1]
      intr_alert_handler_classa, // IDs [145 +: 1]
      intr_otp_ctrl_otp_error, // IDs [144 +: 1]
      intr_otp_ctrl_otp_operation_done, // IDs [143 +: 1]
      1'b0,//intr_usbdev_link_out_err, // IDs [142 +: 1]
      1'b0,//intr_usbdev_connected, // IDs [141 +: 1]
      1'b0,//intr_usbdev_frame, // IDs [140 +: 1]
      1'b0,//intr_usbdev_rx_bitstuff_err, // IDs [139 +: 1]
      1'b0,//intr_usbdev_rx_pid_err, // IDs [138 +: 1]
      1'b0,//1'b0,//intr_usbdev_rx_crc_err, // IDs [137 +: 1]
      1'b0,//intr_usbdev_link_in_err, // IDs [136 +: 1]
      1'b0,//1'b0,//intr_usbdev_av_overflow, // IDs [135 +: 1]
      1'b0,//intr_usbdev_rx_full, // IDs [134 +: 1]
      1'b0,//intr_usbdev_av_empty, // IDs [133 +: 1]
      1'b0,//intr_usbdev_link_resume, // IDs [132 +: 1]
      1'b0,//intr_usbdev_link_suspend, // IDs [131 +: 1]
      1'b0,//intr_usbdev_link_reset, // IDs [130 +: 1]
      1'b0,//intr_usbdev_host_lost, // IDs [129 +: 1]
      1'b0,//intr_usbdev_disconnected, // IDs [128 +: 1]
      1'b0,//intr_usbdev_pkt_sent, // IDs [127 +: 1]
      1'b0,//intr_usbdev_pkt_received, // IDs [126 +: 1]
      intr_rv_timer_timer_expired_0_0, // IDs [125 +: 1]
      1'b0,//intr_pattgen_done_ch1, // IDs [124 +: 1]
      1'b0,//intr_pattgen_done_ch0, // IDs [123 +: 1]
      1'b0,//intr_i2c2_host_timeout, // IDs [122 +: 1]
      1'b0,//intr_i2c2_ack_stop, // IDs [121 +: 1]
      1'b0,//intr_i2c2_acq_overflow, // IDs [120 +: 1]
      1'b0,//intr_i2c2_tx_overflow, // IDs [119 +: 1]
      1'b0,//intr_i2c2_tx_nonempty, // IDs [118 +: 1]
      1'b0,//intr_i2c2_tx_empty, // IDs [117 +: 1]
      1'b0,//intr_i2c2_trans_complete, // IDs [116 +: 1]
      1'b0,//intr_i2c2_sda_unstable, // IDs [115 +: 1]
      1'b0,//intr_i2c2_stretch_timeout, // IDs [114 +: 1]
      1'b0,//intr_i2c2_sda_interference, // IDs [113 +: 1]
      1'b0,//intr_i2c2_scl_interference, // IDs [112 +: 1]
      1'b0,//intr_i2c2_nak, // IDs [111 +: 1]
      1'b0,//intr_i2c2_rx_overflow, // IDs [110 +: 1]
      1'b0,//intr_i2c2_fmt_overflow, // IDs [109 +: 1]
      1'b0,//intr_i2c2_rx_watermark, // IDs [108 +: 1]
      1'b0,//intr_i2c2_fmt_watermark, // IDs [107 +: 1]
      1'b0,//intr_i2c1_host_timeout, // IDs [106 +: 1]
      1'b0,//intr_i2c1_ack_stop, // IDs [105 +: 1]
      1'b0,//intr_i2c1_acq_overflow, // IDs [104 +: 1]
      1'b0,//intr_i2c1_tx_overflow, // IDs [103 +: 1]
      1'b0,//intr_i2c1_tx_nonempty, // IDs [102 +: 1]
      1'b0,//intr_i2c1_tx_empty, // IDs [101 +: 1]
      irq_ibex_i,//1'b0,//intr_i2c1_trans_complete, // IDs [100 +: 1]
      1'b0,//intr_i2c1_sda_unstable, // IDs [99 +: 1]
      1'b0,//intr_i2c1_stretch_timeout, // IDs [98 +: 1]
      1'b0,//intr_i2c1_sda_interference, // IDs [97 +: 1]
      1'b0,//intr_i2c1_scl_interference, // IDs [96 +: 1]
      1'b0,//intr_i2c1_nak, // IDs [95 +: 1]
      1'b0,//intr_i2c1_rx_overflow, // IDs [94 +: 1]
      1'b0,//intr_i2c1_fmt_overflow, // IDs [93 +: 1]
      1'b0,//intr_i2c1_rx_watermark, // IDs [92 +: 1]
      1'b0,//intr_i2c1_fmt_watermark, // IDs [91 +: 1]
      1'b0,//intr_i2c0_host_timeout, // IDs [90 +: 1]
      1'b0,//intr_i2c0_ack_stop, // IDs [89 +: 1]
      1'b0,//intr_i2c0_acq_overflow, // IDs [88 +: 1]
      1'b0,//intr_i2c0_tx_overflow, // IDs [87 +: 1]
      1'b0,//intr_i2c0_tx_nonempty, // IDs [86 +: 1]
      1'b0,//intr_i2c0_tx_empty, // IDs [85 +: 1]
      1'b0,//intr_i2c0_trans_complete, // IDs [84 +: 1]
      1'b0,//intr_i2c0_sda_unstable, // IDs [83 +: 1]
      1'b0,//intr_i2c0_stretch_timeout, // IDs [82 +: 1]
      1'b0,//intr_i2c0_sda_interference, // IDs [81 +: 1]
      1'b0,//intr_i2c0_scl_interference, // IDs [80 +: 1]
      1'b0,//intr_i2c0_nak, // IDs [79 +: 1]
      1'b0,//intr_i2c0_rx_overflow, // IDs [78 +: 1]
      1'b0,//intr_i2c0_fmt_overflow, // IDs [77 +: 1]
      1'b0,//intr_i2c0_rx_watermark, // IDs [76 +: 1]
      1'b0,//intr_i2c0_fmt_watermark, // IDs [75 +: 1]
      1'b0,//intr_spi_host1_spi_event, // IDs [74 +: 1]
      1'b0,//intr_spi_host1_error, // IDs [73 +: 1]
      intr_spi_host0_spi_event, // IDs [72 +: 1]
      intr_spi_host0_error, // IDs [71 +: 1]
      intr_spi_device_txunderflow, // IDs [70 +: 1]
      intr_spi_device_rxoverflow, // IDs [69 +: 1]
      intr_spi_device_rxerr, // IDs [68 +: 1]
      intr_spi_device_txlvl, // IDs [67 +: 1]
      intr_spi_device_rxlvl, // IDs [66 +: 1]
      intr_spi_device_rxf, // IDs [65 +: 1]
      intr_gpio_gpio, // IDs [33 +: 32]
      intr_uart3_rx_parity_err, // IDs [32 +: 1]
      intr_uart3_rx_timeout, // IDs [31 +: 1]
      intr_uart3_rx_break_err, // IDs [30 +: 1]
      intr_uart3_rx_frame_err, // IDs [29 +: 1]
      intr_uart3_rx_overflow, // IDs [28 +: 1]
      intr_uart3_tx_empty, // IDs [27 +: 1]
      intr_uart3_rx_watermark, // IDs [26 +: 1]
      intr_uart3_tx_watermark, // IDs [25 +: 1]
      intr_uart2_rx_parity_err, // IDs [24 +: 1]
      intr_uart2_rx_timeout, // IDs [23 +: 1]
      intr_uart2_rx_break_err, // IDs [22 +: 1]
      intr_uart2_rx_frame_err, // IDs [21 +: 1]
      intr_uart2_rx_overflow, // IDs [20 +: 1]
      intr_uart2_tx_empty, // IDs [19 +: 1]
      intr_uart2_rx_watermark, // IDs [18 +: 1]
      intr_uart2_tx_watermark, // IDs [17 +: 1]
      intr_uart1_rx_parity_err, // IDs [16 +: 1]
      intr_uart1_rx_timeout, // IDs [15 +: 1]
      intr_uart1_rx_break_err, // IDs [14 +: 1]
      intr_uart1_rx_frame_err, // IDs [13 +: 1]
      intr_uart1_rx_overflow, // IDs [12 +: 1]
      intr_uart1_tx_empty, // IDs [11 +: 1]
      intr_uart1_rx_watermark, // IDs [10 +: 1]
      intr_uart1_tx_watermark, // IDs [9 +: 1]
      intr_uart0_rx_parity_err, // IDs [8 +: 1]
      intr_uart0_rx_timeout, // IDs [7 +: 1]
      intr_uart0_rx_break_err, // IDs [6 +: 1]
      intr_uart0_rx_frame_err, // IDs [5 +: 1]
      intr_uart0_rx_overflow, // IDs [4 +: 1]
      intr_uart0_tx_empty, // IDs [3 +: 1]
      intr_uart0_rx_watermark, // IDs [2 +: 1]
      intr_uart0_tx_watermark, // IDs [1 +: 1]
      1'b 0 // ID [0 +: 1] is a special case and tied to zero.
  };

  // TL-UL Crossbar
  xbar_main u_xbar_main (
    .clk_main_i (clkmgr_aon_clocks.clk_main_infra),//clk_main_i),//c
    .clk_fixed_i (clkmgr_aon_clocks.clk_io_div4_infra),//clk_main_i),//
    .rst_main_ni (rstmgr_aon_resets.rst_sys_n[rstmgr_pkg::Domain0Sel]),//por_n_i),//
    .rst_fixed_ni (rstmgr_aon_resets.rst_sys_io_div4_n[rstmgr_pkg::Domain0Sel]),//(por_n_i),//

    // port: tl_rv_core_ibex__corei
    .tl_rv_core_ibex__corei_i(main_tl_rv_core_ibex__corei_req),
    .tl_rv_core_ibex__corei_o(main_tl_rv_core_ibex__corei_rsp),

    // port: tl_rv_core_ibex__cored
    .tl_rv_core_ibex__cored_i(main_tl_rv_core_ibex__cored_req),
    .tl_rv_core_ibex__cored_o(main_tl_rv_core_ibex__cored_rsp),

    //.tl_instr_mem_i(instr2core),
    //.tl_instr_mem_o(core2instr),

    //.tl_ram_2p_i(ram2core),
    //.tl_ram_2p_o(core2ram),

    .tl_sim_ctrl_i(simctrl2core),
    .tl_sim_ctrl_o(core2simctrl),

    .tl_alsaqr_i(alsaqr2core),
    .tl_alsaqr_o(core2alsaqr),

    // port: tl_rv_dm__sba
    .tl_rv_dm__sba_i(main_tl_rv_dm__sba_req),
    .tl_rv_dm__sba_o(main_tl_rv_dm__sba_rsp),

    // port: tl_rv_dm__regs
    .tl_rv_dm__regs_o(rv_dm_regs_tl_d_req),
    .tl_rv_dm__regs_i(rv_dm_regs_tl_d_rsp),

    // port: tl_rv_dm__rom
    .tl_rv_dm__rom_o(rv_dm_rom_tl_d_req),
    .tl_rv_dm__rom_i(rv_dm_rom_tl_d_rsp),

    // port: tl_rom_ctrl__rom
    .tl_rom_ctrl__rom_o(rom_ctrl_rom_tl_req),
    .tl_rom_ctrl__rom_i(rom_ctrl_rom_tl_rsp),

    // port: tl_rom_ctrl__regs
    .tl_rom_ctrl__regs_o(rom_ctrl_regs_tl_req),
    .tl_rom_ctrl__regs_i(rom_ctrl_regs_tl_rsp),

    // port: tl_peri
    .tl_peri_o(main_tl_peri_req),
    .tl_peri_i(main_tl_peri_rsp),

    // port: tl_flash_ctrl__core
    .tl_flash_ctrl__core_o(flash_ctrl_core_tl_req),
    .tl_flash_ctrl__core_i(flash_ctrl_core_tl_rsp),

    // port: tl_flash_ctrl__prim
    .tl_flash_ctrl__prim_o(flash_ctrl_prim_tl_req),
    .tl_flash_ctrl__prim_i(flash_ctrl_prim_tl_rsp),

    // port: tl_flash_ctrl__mem
    .tl_flash_ctrl__mem_o(flash_ctrl_mem_tl_req),
    .tl_flash_ctrl__mem_i(flash_ctrl_mem_tl_rsp),

    // port: tl_hmac
    .tl_hmac_o(hmac_tl_req),
    .tl_hmac_i(hmac_tl_rsp),

    // port: tl_kmac
    .tl_kmac_o(kmac_tl_req),
    .tl_kmac_i(kmac_tl_rsp),

    // port: tl_aes
    .tl_aes_o(aes_tl_req),
    .tl_aes_i(aes_tl_rsp),

    // port: tl_entropy_src
    .tl_entropy_src_o(entropy_src_tl_req),
    .tl_entropy_src_i(entropy_src_tl_rsp),

    // port: tl_csrng
    .tl_csrng_o(csrng_tl_req),
    .tl_csrng_i(csrng_tl_rsp),

    // port: tl_edn0
    .tl_edn0_o(edn0_tl_req),
    .tl_edn0_i(edn0_tl_rsp),

    // port: tl_edn1
    .tl_edn1_o(edn1_tl_req),
    .tl_edn1_i(edn1_tl_rsp),

    // port: tl_rv_plic
    .tl_rv_plic_o(rv_plic_tl_req),
    .tl_rv_plic_i(rv_plic_tl_rsp),

    // port: tl_otbn
    .tl_otbn_o(otbn_tl_req),
    .tl_otbn_i(otbn_tl_rsp),

    // port: tl_keymgr
    .tl_keymgr_o(keymgr_tl_req),
    .tl_keymgr_i(keymgr_tl_rsp),

    // port: tl_rv_core_ibex__cfg
    .tl_rv_core_ibex__cfg_o(rv_core_ibex_cfg_tl_d_req),
    .tl_rv_core_ibex__cfg_i(rv_core_ibex_cfg_tl_d_rsp),

    // port: tl_sram_ctrl_main__regs
    .tl_sram_ctrl_main__regs_o(sram_ctrl_main_regs_tl_req),
    .tl_sram_ctrl_main__regs_i(sram_ctrl_main_regs_tl_rsp),

    // port: tl_sram_ctrl_main__ram
    .tl_sram_ctrl_main__ram_o(sram_ctrl_main_ram_tl_req),//tcore2simctrl),//
    .tl_sram_ctrl_main__ram_i(sram_ctrl_main_ram_tl_rsp),//tsimctrl2core),//

    // port: tl_spi_host0
    .tl_spi_host0_o(spi_host0_tl_req),
    .tl_spi_host0_i(spi_host0_tl_rsp),
/*
    // port: tl_spi_host1
    .tl_spi_host1_o(spi_host1_tl_req),
    .tl_spi_host1_i(spi_host1_tl_rsp),
*/
    .scanmode_i
  );
   
  xbar_peri u_xbar_peri (
    .clk_peri_i (clkmgr_aon_clocks.clk_io_div4_infra),
    .rst_peri_ni (rstmgr_aon_resets.rst_sys_io_div4_n[rstmgr_pkg::Domain0Sel]),

    // port: tl_main
    .tl_main_i(main_tl_peri_req),
    .tl_main_o(main_tl_peri_rsp),

    // port: tl_uart0
    .tl_uart0_o(uart0_tl_req),
    .tl_uart0_i(uart0_tl_rsp),

    // port: tl_uart1
    .tl_uart1_o(uart1_tl_req),
    .tl_uart1_i(uart1_tl_rsp),

    // port: tl_uart2
    .tl_uart2_o(uart2_tl_req),
    .tl_uart2_i(uart2_tl_rsp),

    // port: tl_uart3
    .tl_uart3_o(uart3_tl_req),
    .tl_uart3_i(uart3_tl_rsp),
/*
    // port: tl_i2c0
    .tl_i2c0_o(i2c0_tl_req),
    .tl_i2c0_i(i2c0_tl_rsp),

    // port: tl_i2c1
    .tl_i2c1_o(i2c1_tl_req),
    .tl_i2c1_i(i2c1_tl_rsp),

    // port: tl_i2c2
    .tl_i2c2_o(i2c2_tl_req),
    .tl_i2c2_i(i2c2_tl_rsp),

    // port: tl_pattgen
    .tl_pattgen_o(pattgen_tl_req),
    .tl_pattgen_i(pattgen_tl_rsp),

    // port: tl_pwm_aon
    .tl_pwm_aon_o(pwm_aon_tl_req),
    .tl_pwm_aon_i(pwm_aon_tl_rsp),
*/
    // port: tl_gpio
    .tl_gpio_o(gpio_tl_req),
    .tl_gpio_i(gpio_tl_rsp),

    // port: tl_spi_device
    .tl_spi_device_o(spi_device_tl_req),
    .tl_spi_device_i(spi_device_tl_rsp),

    // port: tl_rv_timer
    .tl_rv_timer_o(rv_timer_tl_req),
    .tl_rv_timer_i(rv_timer_tl_rsp),
/*
    // port: tl_usbdev
    .tl_usbdev_o(usbdev_tl_req),
    .tl_usbdev_i(usbdev_tl_rsp),
*/
    // port: tl_pwrmgr_aon
    .tl_pwrmgr_aon_o(pwrmgr_aon_tl_req),
    .tl_pwrmgr_aon_i(pwrmgr_aon_tl_rsp),

    // port: tl_rstmgr_aon
    .tl_rstmgr_aon_o(rstmgr_aon_tl_req),
    .tl_rstmgr_aon_i(rstmgr_aon_tl_rsp),

    // port: tl_clkmgr_aon
    .tl_clkmgr_aon_o(clkmgr_aon_tl_req),
    .tl_clkmgr_aon_i(clkmgr_aon_tl_rsp),
/*
    // port: tl_pinmux_aon
    .tl_pinmux_aon_o(pinmux_aon_tl_req),
    .tl_pinmux_aon_i(pinmux_aon_tl_rsp),
*/
    // port: tl_otp_ctrl__core
    .tl_otp_ctrl__core_o(otp_ctrl_core_tl_req),
    .tl_otp_ctrl__core_i(otp_ctrl_core_tl_rsp),

    // port: tl_otp_ctrl__prim
    .tl_otp_ctrl__prim_o(otp_ctrl_prim_tl_req),
    .tl_otp_ctrl__prim_i(otp_ctrl_prim_tl_rsp),

    // port: tl_lc_ctrl
    .tl_lc_ctrl_o(lc_ctrl_tl_req),
    .tl_lc_ctrl_i(lc_ctrl_tl_rsp),

    // port: tl_sensor_ctrl_aon
    //.tl_sensor_ctrl_aon_o(sensor_ctrl_aon_tl_req),
    //.tl_sensor_ctrl_aon_i(sensor_ctrl_aon_tl_rsp),

    // port: tl_alert_handler
    .tl_alert_handler_o(alert_handler_tl_req),
    .tl_alert_handler_i(alert_handler_tl_rsp),

    // port: tl_sram_ctrl_ret_aon__regs
    .tl_sram_ctrl_ret_aon__regs_o(sram_ctrl_ret_aon_regs_tl_req),
    .tl_sram_ctrl_ret_aon__regs_i(sram_ctrl_ret_aon_regs_tl_rsp),

    // port: tl_sram_ctrl_ret_aon__ram
    .tl_sram_ctrl_ret_aon__ram_o(sram_ctrl_ret_aon_ram_tl_req),
    .tl_sram_ctrl_ret_aon__ram_i(sram_ctrl_ret_aon_ram_tl_rsp),

    // port: tl_aon_timer_aon
    .tl_aon_timer_aon_o(aon_timer_aon_tl_req),
    .tl_aon_timer_aon_i(aon_timer_aon_tl_rsp),

    // port: tl_sysrst_ctrl_aon
    .tl_sysrst_ctrl_aon_o(sysrst_ctrl_aon_tl_req),
    .tl_sysrst_ctrl_aon_i(sysrst_ctrl_aon_tl_rsp),
/*
    // port: tl_adc_ctrl_aon
    .tl_adc_ctrl_aon_o(adc_ctrl_aon_tl_req),
    .tl_adc_ctrl_aon_i(adc_ctrl_aon_tl_rsp),

    // port: tl_ast
    .tl_ast_o(ast_tl_req_o),
    .tl_ast_i(ast_tl_rsp_i),
*/

    .scanmode_i
  );
  
  // Pinmux connections
  // All muxed inputs
  assign cio_gpio_gpio_p2d[0] = mio_p2d[MioInGpioGpio0];
  assign cio_gpio_gpio_p2d[1] = mio_p2d[MioInGpioGpio1];
  assign cio_gpio_gpio_p2d[2] = mio_p2d[MioInGpioGpio2];
  assign cio_gpio_gpio_p2d[3] = mio_p2d[MioInGpioGpio3];
  assign cio_gpio_gpio_p2d[4] = mio_p2d[MioInGpioGpio4];
  assign cio_gpio_gpio_p2d[5] = mio_p2d[MioInGpioGpio5];
  assign cio_gpio_gpio_p2d[6] = mio_p2d[MioInGpioGpio6];
  assign cio_gpio_gpio_p2d[7] = mio_p2d[MioInGpioGpio7];
  assign cio_gpio_gpio_p2d[8] = mio_p2d[MioInGpioGpio8];
  assign cio_gpio_gpio_p2d[9] = mio_p2d[MioInGpioGpio9];
  assign cio_gpio_gpio_p2d[10] = mio_p2d[MioInGpioGpio10];
  assign cio_gpio_gpio_p2d[11] = mio_p2d[MioInGpioGpio11];
  assign cio_gpio_gpio_p2d[12] = mio_p2d[MioInGpioGpio12];
  assign cio_gpio_gpio_p2d[13] = mio_p2d[MioInGpioGpio13];
  assign cio_gpio_gpio_p2d[14] = mio_p2d[MioInGpioGpio14];
  assign cio_gpio_gpio_p2d[15] = mio_p2d[MioInGpioGpio15];
  assign cio_gpio_gpio_p2d[16] = mio_p2d[MioInGpioGpio16];
  assign cio_gpio_gpio_p2d[17] = mio_p2d[MioInGpioGpio17];
  assign cio_gpio_gpio_p2d[18] = mio_p2d[MioInGpioGpio18];
  assign cio_gpio_gpio_p2d[19] = mio_p2d[MioInGpioGpio19];
  assign cio_gpio_gpio_p2d[20] = mio_p2d[MioInGpioGpio20];
  assign cio_gpio_gpio_p2d[21] = mio_p2d[MioInGpioGpio21];
  assign cio_gpio_gpio_p2d[22] = mio_p2d[MioInGpioGpio22];
  assign cio_gpio_gpio_p2d[23] = mio_p2d[MioInGpioGpio23];
  assign cio_gpio_gpio_p2d[24] = mio_p2d[MioInGpioGpio24];
  assign cio_gpio_gpio_p2d[25] = mio_p2d[MioInGpioGpio25];
  assign cio_gpio_gpio_p2d[26] = mio_p2d[MioInGpioGpio26];
  assign cio_gpio_gpio_p2d[27] = mio_p2d[MioInGpioGpio27];
  assign cio_gpio_gpio_p2d[28] = mio_p2d[MioInGpioGpio28];
  assign cio_gpio_gpio_p2d[29] = mio_p2d[MioInGpioGpio29];
  assign cio_gpio_gpio_p2d[30] = mio_p2d[MioInGpioGpio30];
  assign cio_gpio_gpio_p2d[31] = mio_p2d[MioInGpioGpio31];
  assign cio_i2c0_sda_p2d = mio_p2d[MioInI2c0Sda];
  assign cio_i2c0_scl_p2d = mio_p2d[MioInI2c0Scl];
  assign cio_i2c1_sda_p2d = mio_p2d[MioInI2c1Sda];
  assign cio_i2c1_scl_p2d = mio_p2d[MioInI2c1Scl];
  assign cio_i2c2_sda_p2d = mio_p2d[MioInI2c2Sda];
  assign cio_i2c2_scl_p2d = mio_p2d[MioInI2c2Scl];
  assign cio_spi_host1_sd_p2d[0] = mio_p2d[MioInSpiHost1Sd0];
  assign cio_spi_host1_sd_p2d[1] = mio_p2d[MioInSpiHost1Sd1];
  assign cio_spi_host1_sd_p2d[2] = mio_p2d[MioInSpiHost1Sd2];
  assign cio_spi_host1_sd_p2d[3] = mio_p2d[MioInSpiHost1Sd3];
  assign cio_uart0_rx_p2d = mio_p2d[MioInUart0Rx];
  assign cio_uart1_rx_p2d = mio_p2d[MioInUart1Rx];
  assign cio_uart2_rx_p2d = mio_p2d[MioInUart2Rx];
  assign cio_uart3_rx_p2d = mio_p2d[MioInUart3Rx];
  assign cio_flash_ctrl_tck_p2d = mio_p2d[MioInFlashCtrlTck];
  assign cio_flash_ctrl_tms_p2d = mio_p2d[MioInFlashCtrlTms];
  assign cio_flash_ctrl_tdi_p2d = mio_p2d[MioInFlashCtrlTdi];
  assign cio_sysrst_ctrl_aon_ac_present_p2d = mio_p2d[MioInSysrstCtrlAonAcPresent];
  assign cio_sysrst_ctrl_aon_key0_in_p2d = 1'b0;//mio_p2d[MioInSysrstCtrlAonKey0In];
  assign cio_sysrst_ctrl_aon_key1_in_p2d = 1'b0;//mio_p2d[MioInSysrstCtrlAonKey1In];
  assign cio_sysrst_ctrl_aon_key2_in_p2d = 1'b0;//mio_p2d[MioInSysrstCtrlAonKey2In];
  assign cio_sysrst_ctrl_aon_pwrb_in_p2d = 1'b0;//mio_p2d[MioInSysrstCtrlAonPwrbIn];
  assign cio_sysrst_ctrl_aon_lid_open_p2d = mio_p2d[MioInSysrstCtrlAonLidOpen];

  // All muxed outputs
  assign mio_d2p[MioOutGpioGpio0] = cio_gpio_gpio_d2p[0];
  assign mio_d2p[MioOutGpioGpio1] = cio_gpio_gpio_d2p[1];
  assign mio_d2p[MioOutGpioGpio2] = cio_gpio_gpio_d2p[2];
  assign mio_d2p[MioOutGpioGpio3] = cio_gpio_gpio_d2p[3];
  assign mio_d2p[MioOutGpioGpio4] = cio_gpio_gpio_d2p[4];
  assign mio_d2p[MioOutGpioGpio5] = cio_gpio_gpio_d2p[5];
  assign mio_d2p[MioOutGpioGpio6] = cio_gpio_gpio_d2p[6];
  assign mio_d2p[MioOutGpioGpio7] = cio_gpio_gpio_d2p[7];
  assign mio_d2p[MioOutGpioGpio8] = cio_gpio_gpio_d2p[8];
  assign mio_d2p[MioOutGpioGpio9] = cio_gpio_gpio_d2p[9];
  assign mio_d2p[MioOutGpioGpio10] = cio_gpio_gpio_d2p[10];
  assign mio_d2p[MioOutGpioGpio11] = cio_gpio_gpio_d2p[11];
  assign mio_d2p[MioOutGpioGpio12] = cio_gpio_gpio_d2p[12];
  assign mio_d2p[MioOutGpioGpio13] = cio_gpio_gpio_d2p[13];
  assign mio_d2p[MioOutGpioGpio14] = cio_gpio_gpio_d2p[14];
  assign mio_d2p[MioOutGpioGpio15] = cio_gpio_gpio_d2p[15];
  assign mio_d2p[MioOutGpioGpio16] = cio_gpio_gpio_d2p[16];
  assign mio_d2p[MioOutGpioGpio17] = cio_gpio_gpio_d2p[17];
  assign mio_d2p[MioOutGpioGpio18] = cio_gpio_gpio_d2p[18];
  assign mio_d2p[MioOutGpioGpio19] = cio_gpio_gpio_d2p[19];
  assign mio_d2p[MioOutGpioGpio20] = cio_gpio_gpio_d2p[20];
  assign mio_d2p[MioOutGpioGpio21] = cio_gpio_gpio_d2p[21];
  assign mio_d2p[MioOutGpioGpio22] = cio_gpio_gpio_d2p[22];
  assign mio_d2p[MioOutGpioGpio23] = cio_gpio_gpio_d2p[23];
  assign mio_d2p[MioOutGpioGpio24] = cio_gpio_gpio_d2p[24];
  assign mio_d2p[MioOutGpioGpio25] = cio_gpio_gpio_d2p[25];
  assign mio_d2p[MioOutGpioGpio26] = cio_gpio_gpio_d2p[26];
  assign mio_d2p[MioOutGpioGpio27] = cio_gpio_gpio_d2p[27];
  assign mio_d2p[MioOutGpioGpio28] = cio_gpio_gpio_d2p[28];
  assign mio_d2p[MioOutGpioGpio29] = cio_gpio_gpio_d2p[29];
  assign mio_d2p[MioOutGpioGpio30] = cio_gpio_gpio_d2p[30];
  assign mio_d2p[MioOutGpioGpio31] = cio_gpio_gpio_d2p[31];
  assign mio_d2p[MioOutI2c0Sda] = cio_i2c0_sda_d2p;
  assign mio_d2p[MioOutI2c0Scl] = cio_i2c0_scl_d2p;
  assign mio_d2p[MioOutI2c1Sda] = cio_i2c1_sda_d2p;
  assign mio_d2p[MioOutI2c1Scl] = cio_i2c1_scl_d2p;
  assign mio_d2p[MioOutI2c2Sda] = cio_i2c2_sda_d2p;
  assign mio_d2p[MioOutI2c2Scl] = cio_i2c2_scl_d2p;
  assign mio_d2p[MioOutSpiHost1Sd0] = cio_spi_host1_sd_d2p[0];
  assign mio_d2p[MioOutSpiHost1Sd1] = cio_spi_host1_sd_d2p[1];
  assign mio_d2p[MioOutSpiHost1Sd2] = cio_spi_host1_sd_d2p[2];
  assign mio_d2p[MioOutSpiHost1Sd3] = cio_spi_host1_sd_d2p[3];
  assign mio_d2p[MioOutUart0Tx] = cio_uart0_tx_d2p;
  assign mio_d2p[MioOutUart1Tx] = cio_uart1_tx_d2p;
  assign mio_d2p[MioOutUart2Tx] = cio_uart2_tx_d2p;
  assign mio_d2p[MioOutUart3Tx] = cio_uart3_tx_d2p;
  assign mio_d2p[MioOutPattgenPda0Tx] = cio_pattgen_pda0_tx_d2p;
  assign mio_d2p[MioOutPattgenPcl0Tx] = cio_pattgen_pcl0_tx_d2p;
  assign mio_d2p[MioOutPattgenPda1Tx] = cio_pattgen_pda1_tx_d2p;
  assign mio_d2p[MioOutPattgenPcl1Tx] = cio_pattgen_pcl1_tx_d2p;
  assign mio_d2p[MioOutSpiHost1Sck] = cio_spi_host1_sck_d2p;
  assign mio_d2p[MioOutSpiHost1Csb] = cio_spi_host1_csb_d2p;
  assign mio_d2p[MioOutFlashCtrlTdo] = cio_flash_ctrl_tdo_d2p;
  assign mio_d2p[MioOutSensorCtrlAonAstDebugOut0] = cio_sensor_ctrl_aon_ast_debug_out_d2p[0];
  assign mio_d2p[MioOutSensorCtrlAonAstDebugOut1] = cio_sensor_ctrl_aon_ast_debug_out_d2p[1];
  assign mio_d2p[MioOutSensorCtrlAonAstDebugOut2] = cio_sensor_ctrl_aon_ast_debug_out_d2p[2];
  assign mio_d2p[MioOutSensorCtrlAonAstDebugOut3] = cio_sensor_ctrl_aon_ast_debug_out_d2p[3];
  assign mio_d2p[MioOutSensorCtrlAonAstDebugOut4] = cio_sensor_ctrl_aon_ast_debug_out_d2p[4];
  assign mio_d2p[MioOutSensorCtrlAonAstDebugOut5] = cio_sensor_ctrl_aon_ast_debug_out_d2p[5];
  assign mio_d2p[MioOutSensorCtrlAonAstDebugOut6] = cio_sensor_ctrl_aon_ast_debug_out_d2p[6];
  assign mio_d2p[MioOutSensorCtrlAonAstDebugOut7] = cio_sensor_ctrl_aon_ast_debug_out_d2p[7];
  assign mio_d2p[MioOutSensorCtrlAonAstDebugOut8] = cio_sensor_ctrl_aon_ast_debug_out_d2p[8];
  assign mio_d2p[MioOutPwmAonPwm0] = cio_pwm_aon_pwm_d2p[0];
  assign mio_d2p[MioOutPwmAonPwm1] = cio_pwm_aon_pwm_d2p[1];
  assign mio_d2p[MioOutPwmAonPwm2] = cio_pwm_aon_pwm_d2p[2];
  assign mio_d2p[MioOutPwmAonPwm3] = cio_pwm_aon_pwm_d2p[3];
  assign mio_d2p[MioOutPwmAonPwm4] = cio_pwm_aon_pwm_d2p[4];
  assign mio_d2p[MioOutPwmAonPwm5] = cio_pwm_aon_pwm_d2p[5];
  assign mio_d2p[MioOutOtpCtrlTest0] = cio_otp_ctrl_test_d2p[0];
  assign mio_d2p[MioOutSysrstCtrlAonBatDisable] = cio_sysrst_ctrl_aon_bat_disable_d2p;
  assign mio_d2p[MioOutSysrstCtrlAonKey0Out] = cio_sysrst_ctrl_aon_key0_out_d2p;
  assign mio_d2p[MioOutSysrstCtrlAonKey1Out] = cio_sysrst_ctrl_aon_key1_out_d2p;
  assign mio_d2p[MioOutSysrstCtrlAonKey2Out] = cio_sysrst_ctrl_aon_key2_out_d2p;
  assign mio_d2p[MioOutSysrstCtrlAonPwrbOut] = cio_sysrst_ctrl_aon_pwrb_out_d2p;
  assign mio_d2p[MioOutSysrstCtrlAonZ3Wakeup] = cio_sysrst_ctrl_aon_z3_wakeup_d2p;

  // All muxed output enables
  assign mio_en_d2p[MioOutGpioGpio0] = cio_gpio_gpio_en_d2p[0];
  assign mio_en_d2p[MioOutGpioGpio1] = cio_gpio_gpio_en_d2p[1];
  assign mio_en_d2p[MioOutGpioGpio2] = cio_gpio_gpio_en_d2p[2];
  assign mio_en_d2p[MioOutGpioGpio3] = cio_gpio_gpio_en_d2p[3];
  assign mio_en_d2p[MioOutGpioGpio4] = cio_gpio_gpio_en_d2p[4];
  assign mio_en_d2p[MioOutGpioGpio5] = cio_gpio_gpio_en_d2p[5];
  assign mio_en_d2p[MioOutGpioGpio6] = cio_gpio_gpio_en_d2p[6];
  assign mio_en_d2p[MioOutGpioGpio7] = cio_gpio_gpio_en_d2p[7];
  assign mio_en_d2p[MioOutGpioGpio8] = cio_gpio_gpio_en_d2p[8];
  assign mio_en_d2p[MioOutGpioGpio9] = cio_gpio_gpio_en_d2p[9];
  assign mio_en_d2p[MioOutGpioGpio10] = cio_gpio_gpio_en_d2p[10];
  assign mio_en_d2p[MioOutGpioGpio11] = cio_gpio_gpio_en_d2p[11];
  assign mio_en_d2p[MioOutGpioGpio12] = cio_gpio_gpio_en_d2p[12];
  assign mio_en_d2p[MioOutGpioGpio13] = cio_gpio_gpio_en_d2p[13];
  assign mio_en_d2p[MioOutGpioGpio14] = cio_gpio_gpio_en_d2p[14];
  assign mio_en_d2p[MioOutGpioGpio15] = cio_gpio_gpio_en_d2p[15];
  assign mio_en_d2p[MioOutGpioGpio16] = cio_gpio_gpio_en_d2p[16];
  assign mio_en_d2p[MioOutGpioGpio17] = cio_gpio_gpio_en_d2p[17];
  assign mio_en_d2p[MioOutGpioGpio18] = cio_gpio_gpio_en_d2p[18];
  assign mio_en_d2p[MioOutGpioGpio19] = cio_gpio_gpio_en_d2p[19];
  assign mio_en_d2p[MioOutGpioGpio20] = cio_gpio_gpio_en_d2p[20];
  assign mio_en_d2p[MioOutGpioGpio21] = cio_gpio_gpio_en_d2p[21];
  assign mio_en_d2p[MioOutGpioGpio22] = cio_gpio_gpio_en_d2p[22];
  assign mio_en_d2p[MioOutGpioGpio23] = cio_gpio_gpio_en_d2p[23];
  assign mio_en_d2p[MioOutGpioGpio24] = cio_gpio_gpio_en_d2p[24];
  assign mio_en_d2p[MioOutGpioGpio25] = cio_gpio_gpio_en_d2p[25];
  assign mio_en_d2p[MioOutGpioGpio26] = cio_gpio_gpio_en_d2p[26];
  assign mio_en_d2p[MioOutGpioGpio27] = cio_gpio_gpio_en_d2p[27];
  assign mio_en_d2p[MioOutGpioGpio28] = cio_gpio_gpio_en_d2p[28];
  assign mio_en_d2p[MioOutGpioGpio29] = cio_gpio_gpio_en_d2p[29];
  assign mio_en_d2p[MioOutGpioGpio30] = cio_gpio_gpio_en_d2p[30];
  assign mio_en_d2p[MioOutGpioGpio31] = cio_gpio_gpio_en_d2p[31];
  assign mio_en_d2p[MioOutI2c0Sda] = cio_i2c0_sda_en_d2p;
  assign mio_en_d2p[MioOutI2c0Scl] = cio_i2c0_scl_en_d2p;
  assign mio_en_d2p[MioOutI2c1Sda] = cio_i2c1_sda_en_d2p;
  assign mio_en_d2p[MioOutI2c1Scl] = cio_i2c1_scl_en_d2p;
  assign mio_en_d2p[MioOutI2c2Sda] = cio_i2c2_sda_en_d2p;
  assign mio_en_d2p[MioOutI2c2Scl] = cio_i2c2_scl_en_d2p;
  assign mio_en_d2p[MioOutSpiHost1Sd0] = cio_spi_host1_sd_en_d2p[0];
  assign mio_en_d2p[MioOutSpiHost1Sd1] = cio_spi_host1_sd_en_d2p[1];
  assign mio_en_d2p[MioOutSpiHost1Sd2] = cio_spi_host1_sd_en_d2p[2];
  assign mio_en_d2p[MioOutSpiHost1Sd3] = cio_spi_host1_sd_en_d2p[3];
  assign mio_en_d2p[MioOutUart0Tx] = cio_uart0_tx_en_d2p;
  assign mio_en_d2p[MioOutUart1Tx] = cio_uart1_tx_en_d2p;
  assign mio_en_d2p[MioOutUart2Tx] = cio_uart2_tx_en_d2p;
  assign mio_en_d2p[MioOutUart3Tx] = cio_uart3_tx_en_d2p;
  assign mio_en_d2p[MioOutPattgenPda0Tx] = cio_pattgen_pda0_tx_en_d2p;
  assign mio_en_d2p[MioOutPattgenPcl0Tx] = cio_pattgen_pcl0_tx_en_d2p;
  assign mio_en_d2p[MioOutPattgenPda1Tx] = cio_pattgen_pda1_tx_en_d2p;
  assign mio_en_d2p[MioOutPattgenPcl1Tx] = cio_pattgen_pcl1_tx_en_d2p;
  assign mio_en_d2p[MioOutSpiHost1Sck] = cio_spi_host1_sck_en_d2p;
  assign mio_en_d2p[MioOutSpiHost1Csb] = cio_spi_host1_csb_en_d2p;
  assign mio_en_d2p[MioOutFlashCtrlTdo] = cio_flash_ctrl_tdo_en_d2p;
  assign mio_en_d2p[MioOutSensorCtrlAonAstDebugOut0] = cio_sensor_ctrl_aon_ast_debug_out_en_d2p[0];
  assign mio_en_d2p[MioOutSensorCtrlAonAstDebugOut1] = cio_sensor_ctrl_aon_ast_debug_out_en_d2p[1];
  assign mio_en_d2p[MioOutSensorCtrlAonAstDebugOut2] = cio_sensor_ctrl_aon_ast_debug_out_en_d2p[2];
  assign mio_en_d2p[MioOutSensorCtrlAonAstDebugOut3] = cio_sensor_ctrl_aon_ast_debug_out_en_d2p[3];
  assign mio_en_d2p[MioOutSensorCtrlAonAstDebugOut4] = cio_sensor_ctrl_aon_ast_debug_out_en_d2p[4];
  assign mio_en_d2p[MioOutSensorCtrlAonAstDebugOut5] = cio_sensor_ctrl_aon_ast_debug_out_en_d2p[5];
  assign mio_en_d2p[MioOutSensorCtrlAonAstDebugOut6] = cio_sensor_ctrl_aon_ast_debug_out_en_d2p[6];
  assign mio_en_d2p[MioOutSensorCtrlAonAstDebugOut7] = cio_sensor_ctrl_aon_ast_debug_out_en_d2p[7];
  assign mio_en_d2p[MioOutSensorCtrlAonAstDebugOut8] = cio_sensor_ctrl_aon_ast_debug_out_en_d2p[8];
  assign mio_en_d2p[MioOutPwmAonPwm0] = cio_pwm_aon_pwm_en_d2p[0];
  assign mio_en_d2p[MioOutPwmAonPwm1] = cio_pwm_aon_pwm_en_d2p[1];
  assign mio_en_d2p[MioOutPwmAonPwm2] = cio_pwm_aon_pwm_en_d2p[2];
  assign mio_en_d2p[MioOutPwmAonPwm3] = cio_pwm_aon_pwm_en_d2p[3];
  assign mio_en_d2p[MioOutPwmAonPwm4] = cio_pwm_aon_pwm_en_d2p[4];
  assign mio_en_d2p[MioOutPwmAonPwm5] = cio_pwm_aon_pwm_en_d2p[5];
  assign mio_en_d2p[MioOutOtpCtrlTest0] = cio_otp_ctrl_test_en_d2p[0];
  assign mio_en_d2p[MioOutSysrstCtrlAonBatDisable] = cio_sysrst_ctrl_aon_bat_disable_en_d2p;
  assign mio_en_d2p[MioOutSysrstCtrlAonKey0Out] = cio_sysrst_ctrl_aon_key0_out_en_d2p;
  assign mio_en_d2p[MioOutSysrstCtrlAonKey1Out] = cio_sysrst_ctrl_aon_key1_out_en_d2p;
  assign mio_en_d2p[MioOutSysrstCtrlAonKey2Out] = cio_sysrst_ctrl_aon_key2_out_en_d2p;
  assign mio_en_d2p[MioOutSysrstCtrlAonPwrbOut] = cio_sysrst_ctrl_aon_pwrb_out_en_d2p;
  assign mio_en_d2p[MioOutSysrstCtrlAonZ3Wakeup] = cio_sysrst_ctrl_aon_z3_wakeup_en_d2p;

  // All dedicated inputs
  logic [23:0] unused_dio_p2d;
  assign unused_dio_p2d = dio_p2d;
 
  assign cio_usbdev_d_p2d = dio_p2d[DioUsbdevD];
  assign cio_usbdev_dp_p2d = dio_p2d[DioUsbdevDp];
  assign cio_usbdev_dn_p2d = dio_p2d[DioUsbdevDn];
  assign cio_sysrst_ctrl_aon_ec_rst_l_p2d = dio_p2d[DioSysrstCtrlAonEcRstL];
  assign cio_usbdev_sense_p2d = dio_p2d[DioUsbdevSense];

    // All dedicated outputs
  assign dio_d2p[DioSpiHost0Sd0] = cio_spi_host0_sd_d2p[0];
  assign dio_d2p[DioSpiHost0Sd1] = cio_spi_host0_sd_d2p[1];
  assign dio_d2p[DioSpiHost0Sd2] = cio_spi_host0_sd_d2p[2];
  assign dio_d2p[DioSpiHost0Sd3] = cio_spi_host0_sd_d2p[3];
  assign dio_d2p[DioSpiDeviceSd0] = cio_spi_device_sd_d2p[0];
  assign dio_d2p[DioSpiDeviceSd1] = cio_spi_device_sd_d2p[1];
  assign dio_d2p[DioSpiDeviceSd2] = cio_spi_device_sd_d2p[2];
  assign dio_d2p[DioSpiDeviceSd3] = cio_spi_device_sd_d2p[3];
  assign dio_d2p[DioUsbdevD] = cio_usbdev_d_d2p;
  assign dio_d2p[DioUsbdevDp] = cio_usbdev_dp_d2p;
  assign dio_d2p[DioUsbdevDn] = cio_usbdev_dn_d2p;
  assign dio_d2p[DioSysrstCtrlAonEcRstL] = cio_sysrst_ctrl_aon_ec_rst_l_d2p;
  assign dio_d2p[DioSpiDeviceSck] = 1'b0;
  assign dio_d2p[DioSpiDeviceCsb] = 1'b0;
  assign dio_d2p[DioUsbdevSense] = 1'b0;
  assign dio_d2p[DioSpiHost0Sck] = cio_spi_host0_sck_d2p;
  assign dio_d2p[DioSpiHost0Csb] = cio_spi_host0_csb_d2p;
  assign dio_d2p[DioUsbdevSe0] = cio_usbdev_se0_d2p;
  assign dio_d2p[DioUsbdevDpPullup] = cio_usbdev_dp_pullup_d2p;
  assign dio_d2p[DioUsbdevDnPullup] = cio_usbdev_dn_pullup_d2p;
  assign dio_d2p[DioUsbdevTxModeSe] = cio_usbdev_tx_mode_se_d2p;
  assign dio_d2p[DioUsbdevSuspend] = cio_usbdev_suspend_d2p;
  assign dio_d2p[DioUsbdevRxEnable] = cio_usbdev_rx_enable_d2p;
  assign dio_d2p[DioSysrstCtrlAonFlashWpL] = cio_sysrst_ctrl_aon_flash_wp_l_d2p;

  // All dedicated output enables
  assign dio_en_d2p[DioSpiHost0Sd0] = cio_spi_host0_sd_en_d2p[0];
  assign dio_en_d2p[DioSpiHost0Sd1] = cio_spi_host0_sd_en_d2p[1];
  assign dio_en_d2p[DioSpiHost0Sd2] = cio_spi_host0_sd_en_d2p[2];
  assign dio_en_d2p[DioSpiHost0Sd3] = cio_spi_host0_sd_en_d2p[3];
  assign dio_en_d2p[DioSpiDeviceSd0] = cio_spi_device_sd_en_d2p[0];
  assign dio_en_d2p[DioSpiDeviceSd1] = cio_spi_device_sd_en_d2p[1];
  assign dio_en_d2p[DioSpiDeviceSd2] = cio_spi_device_sd_en_d2p[2];
  assign dio_en_d2p[DioSpiDeviceSd3] = cio_spi_device_sd_en_d2p[3];
  assign dio_en_d2p[DioUsbdevD] = cio_usbdev_d_en_d2p;
  assign dio_en_d2p[DioUsbdevDp] = cio_usbdev_dp_en_d2p;
  assign dio_en_d2p[DioUsbdevDn] = cio_usbdev_dn_en_d2p;
  assign dio_en_d2p[DioSysrstCtrlAonEcRstL] = cio_sysrst_ctrl_aon_ec_rst_l_en_d2p;
  assign dio_en_d2p[DioSpiDeviceSck] = 1'b0;
  assign dio_en_d2p[DioSpiDeviceCsb] = 1'b0;
  assign dio_en_d2p[DioUsbdevSense] = 1'b0;
  assign dio_en_d2p[DioSpiHost0Sck] = cio_spi_host0_sck_en_d2p;
  assign dio_en_d2p[DioSpiHost0Csb] = cio_spi_host0_csb_en_d2p;
  assign dio_en_d2p[DioUsbdevSe0] = cio_usbdev_se0_en_d2p;
  assign dio_en_d2p[DioUsbdevDpPullup] = cio_usbdev_dp_pullup_en_d2p;
  assign dio_en_d2p[DioUsbdevDnPullup] = cio_usbdev_dn_pullup_en_d2p;
  assign dio_en_d2p[DioUsbdevTxModeSe] = cio_usbdev_tx_mode_se_en_d2p;
  assign dio_en_d2p[DioUsbdevSuspend] = cio_usbdev_suspend_en_d2p;
  assign dio_en_d2p[DioUsbdevRxEnable] = cio_usbdev_rx_enable_en_d2p;
  assign dio_en_d2p[DioSysrstCtrlAonFlashWpL] = cio_sysrst_ctrl_aon_flash_wp_l_en_d2p;


  // make sure scanmode_i is never X (including during reset)
  `ASSERT_KNOWN(scanmodeKnown, scanmode_i, clk_main_i, 0)


endmodule
